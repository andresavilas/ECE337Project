library verilog;
use verilog.vl_types.all;
entity tb_miner_core_sma is
end tb_miner_core_sma;
