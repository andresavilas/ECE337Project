library verilog;
use verilog.vl_types.all;
entity tb_miner_core_sha is
end tb_miner_core_sha;
