
module uart_tx_TCU ( clk, n_rst, send_data, done, tim_en, load_en );
  input clk, n_rst, send_data, done;
  output tim_en, load_en;
  wire   state, n5, n2, n3;
  assign tim_en = state;

  DFFSR state_reg ( .D(n5), .CLK(clk), .R(n_rst), .S(1'b1), .Q(state) );
  INVX1 U3 ( .A(n2), .Y(load_en) );
  OAI21X1 U4 ( .A(done), .B(n3), .C(n2), .Y(n5) );
  NAND2X1 U5 ( .A(send_data), .B(n3), .Y(n2) );
  INVX1 U6 ( .A(state), .Y(n3) );
endmodule


module flex_pts_sr_NUM_BITS360_SHIFT_MSB1 ( clk, n_rst, shift_enable, 
        load_enable, parallel_in, serial_out );
  input [359:0] parallel_in;
  input clk, n_rst, shift_enable, load_enable;
  output serial_out;
  wire   n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557;
  wire   [358:0] buffer;

  DFFSR \buffer_reg[0]  ( .D(n1444), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[0]) );
  DFFSR \buffer_reg[1]  ( .D(n1443), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[1]) );
  DFFSR \buffer_reg[2]  ( .D(n1442), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[2]) );
  DFFSR \buffer_reg[3]  ( .D(n1441), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[3]) );
  DFFSR \buffer_reg[4]  ( .D(n1440), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[4]) );
  DFFSR \buffer_reg[5]  ( .D(n1439), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[5]) );
  DFFSR \buffer_reg[6]  ( .D(n1438), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[6]) );
  DFFSR \buffer_reg[7]  ( .D(n1437), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[7]) );
  DFFSR \buffer_reg[8]  ( .D(n1436), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[8]) );
  DFFSR \buffer_reg[9]  ( .D(n1435), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[9]) );
  DFFSR \buffer_reg[10]  ( .D(n1434), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[10]) );
  DFFSR \buffer_reg[11]  ( .D(n1433), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[11]) );
  DFFSR \buffer_reg[12]  ( .D(n1432), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[12]) );
  DFFSR \buffer_reg[13]  ( .D(n1431), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[13]) );
  DFFSR \buffer_reg[14]  ( .D(n1430), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[14]) );
  DFFSR \buffer_reg[15]  ( .D(n1429), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[15]) );
  DFFSR \buffer_reg[16]  ( .D(n1428), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[16]) );
  DFFSR \buffer_reg[17]  ( .D(n1427), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[17]) );
  DFFSR \buffer_reg[18]  ( .D(n1426), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[18]) );
  DFFSR \buffer_reg[19]  ( .D(n1425), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[19]) );
  DFFSR \buffer_reg[20]  ( .D(n1424), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[20]) );
  DFFSR \buffer_reg[21]  ( .D(n1423), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[21]) );
  DFFSR \buffer_reg[22]  ( .D(n1422), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[22]) );
  DFFSR \buffer_reg[23]  ( .D(n1421), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[23]) );
  DFFSR \buffer_reg[24]  ( .D(n1420), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[24]) );
  DFFSR \buffer_reg[25]  ( .D(n1419), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[25]) );
  DFFSR \buffer_reg[26]  ( .D(n1418), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[26]) );
  DFFSR \buffer_reg[27]  ( .D(n1417), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[27]) );
  DFFSR \buffer_reg[28]  ( .D(n1416), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[28]) );
  DFFSR \buffer_reg[29]  ( .D(n1415), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[29]) );
  DFFSR \buffer_reg[30]  ( .D(n1414), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[30]) );
  DFFSR \buffer_reg[31]  ( .D(n1413), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[31]) );
  DFFSR \buffer_reg[32]  ( .D(n1412), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[32]) );
  DFFSR \buffer_reg[33]  ( .D(n1411), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[33]) );
  DFFSR \buffer_reg[34]  ( .D(n1410), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[34]) );
  DFFSR \buffer_reg[35]  ( .D(n1409), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[35]) );
  DFFSR \buffer_reg[36]  ( .D(n1408), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[36]) );
  DFFSR \buffer_reg[37]  ( .D(n1407), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[37]) );
  DFFSR \buffer_reg[38]  ( .D(n1406), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[38]) );
  DFFSR \buffer_reg[39]  ( .D(n1405), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[39]) );
  DFFSR \buffer_reg[40]  ( .D(n1404), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[40]) );
  DFFSR \buffer_reg[41]  ( .D(n1403), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[41]) );
  DFFSR \buffer_reg[42]  ( .D(n1402), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[42]) );
  DFFSR \buffer_reg[43]  ( .D(n1401), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[43]) );
  DFFSR \buffer_reg[44]  ( .D(n1400), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[44]) );
  DFFSR \buffer_reg[45]  ( .D(n1399), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[45]) );
  DFFSR \buffer_reg[46]  ( .D(n1398), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[46]) );
  DFFSR \buffer_reg[47]  ( .D(n1397), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[47]) );
  DFFSR \buffer_reg[48]  ( .D(n1396), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[48]) );
  DFFSR \buffer_reg[49]  ( .D(n1395), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[49]) );
  DFFSR \buffer_reg[50]  ( .D(n1394), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[50]) );
  DFFSR \buffer_reg[51]  ( .D(n1393), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[51]) );
  DFFSR \buffer_reg[52]  ( .D(n1392), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[52]) );
  DFFSR \buffer_reg[53]  ( .D(n1391), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[53]) );
  DFFSR \buffer_reg[54]  ( .D(n1390), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[54]) );
  DFFSR \buffer_reg[55]  ( .D(n1389), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[55]) );
  DFFSR \buffer_reg[56]  ( .D(n1388), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[56]) );
  DFFSR \buffer_reg[57]  ( .D(n1387), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[57]) );
  DFFSR \buffer_reg[58]  ( .D(n1386), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[58]) );
  DFFSR \buffer_reg[59]  ( .D(n1385), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[59]) );
  DFFSR \buffer_reg[60]  ( .D(n1384), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[60]) );
  DFFSR \buffer_reg[61]  ( .D(n1383), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[61]) );
  DFFSR \buffer_reg[62]  ( .D(n1382), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[62]) );
  DFFSR \buffer_reg[63]  ( .D(n1381), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[63]) );
  DFFSR \buffer_reg[64]  ( .D(n1380), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[64]) );
  DFFSR \buffer_reg[65]  ( .D(n1379), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[65]) );
  DFFSR \buffer_reg[66]  ( .D(n1378), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[66]) );
  DFFSR \buffer_reg[67]  ( .D(n1377), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[67]) );
  DFFSR \buffer_reg[68]  ( .D(n1376), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[68]) );
  DFFSR \buffer_reg[69]  ( .D(n1375), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[69]) );
  DFFSR \buffer_reg[70]  ( .D(n1374), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[70]) );
  DFFSR \buffer_reg[71]  ( .D(n1373), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[71]) );
  DFFSR \buffer_reg[72]  ( .D(n1372), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[72]) );
  DFFSR \buffer_reg[73]  ( .D(n1371), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[73]) );
  DFFSR \buffer_reg[74]  ( .D(n1370), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[74]) );
  DFFSR \buffer_reg[75]  ( .D(n1369), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[75]) );
  DFFSR \buffer_reg[76]  ( .D(n1368), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[76]) );
  DFFSR \buffer_reg[77]  ( .D(n1367), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[77]) );
  DFFSR \buffer_reg[78]  ( .D(n1366), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[78]) );
  DFFSR \buffer_reg[79]  ( .D(n1365), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[79]) );
  DFFSR \buffer_reg[80]  ( .D(n1364), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[80]) );
  DFFSR \buffer_reg[81]  ( .D(n1363), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[81]) );
  DFFSR \buffer_reg[82]  ( .D(n1362), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[82]) );
  DFFSR \buffer_reg[83]  ( .D(n1361), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[83]) );
  DFFSR \buffer_reg[84]  ( .D(n1360), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[84]) );
  DFFSR \buffer_reg[85]  ( .D(n1359), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[85]) );
  DFFSR \buffer_reg[86]  ( .D(n1358), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[86]) );
  DFFSR \buffer_reg[87]  ( .D(n1357), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[87]) );
  DFFSR \buffer_reg[88]  ( .D(n1356), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[88]) );
  DFFSR \buffer_reg[89]  ( .D(n1355), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[89]) );
  DFFSR \buffer_reg[90]  ( .D(n1354), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[90]) );
  DFFSR \buffer_reg[91]  ( .D(n1353), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[91]) );
  DFFSR \buffer_reg[92]  ( .D(n1352), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[92]) );
  DFFSR \buffer_reg[93]  ( .D(n1351), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[93]) );
  DFFSR \buffer_reg[94]  ( .D(n1350), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[94]) );
  DFFSR \buffer_reg[95]  ( .D(n1349), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[95]) );
  DFFSR \buffer_reg[96]  ( .D(n1348), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[96]) );
  DFFSR \buffer_reg[97]  ( .D(n1347), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[97]) );
  DFFSR \buffer_reg[98]  ( .D(n1346), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[98]) );
  DFFSR \buffer_reg[99]  ( .D(n1345), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[99]) );
  DFFSR \buffer_reg[100]  ( .D(n1344), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[100]) );
  DFFSR \buffer_reg[101]  ( .D(n1343), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[101]) );
  DFFSR \buffer_reg[102]  ( .D(n1342), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[102]) );
  DFFSR \buffer_reg[103]  ( .D(n1341), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[103]) );
  DFFSR \buffer_reg[104]  ( .D(n1340), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[104]) );
  DFFSR \buffer_reg[105]  ( .D(n1339), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[105]) );
  DFFSR \buffer_reg[106]  ( .D(n1338), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[106]) );
  DFFSR \buffer_reg[107]  ( .D(n1337), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[107]) );
  DFFSR \buffer_reg[108]  ( .D(n1336), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[108]) );
  DFFSR \buffer_reg[109]  ( .D(n1335), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[109]) );
  DFFSR \buffer_reg[110]  ( .D(n1334), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[110]) );
  DFFSR \buffer_reg[111]  ( .D(n1333), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[111]) );
  DFFSR \buffer_reg[112]  ( .D(n1332), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[112]) );
  DFFSR \buffer_reg[113]  ( .D(n1331), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[113]) );
  DFFSR \buffer_reg[114]  ( .D(n1330), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[114]) );
  DFFSR \buffer_reg[115]  ( .D(n1329), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[115]) );
  DFFSR \buffer_reg[116]  ( .D(n1328), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[116]) );
  DFFSR \buffer_reg[117]  ( .D(n1327), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[117]) );
  DFFSR \buffer_reg[118]  ( .D(n1326), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[118]) );
  DFFSR \buffer_reg[119]  ( .D(n1325), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[119]) );
  DFFSR \buffer_reg[120]  ( .D(n1324), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[120]) );
  DFFSR \buffer_reg[121]  ( .D(n1323), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[121]) );
  DFFSR \buffer_reg[122]  ( .D(n1322), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[122]) );
  DFFSR \buffer_reg[123]  ( .D(n1321), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[123]) );
  DFFSR \buffer_reg[124]  ( .D(n1320), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[124]) );
  DFFSR \buffer_reg[125]  ( .D(n1319), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[125]) );
  DFFSR \buffer_reg[126]  ( .D(n1318), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[126]) );
  DFFSR \buffer_reg[127]  ( .D(n1317), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[127]) );
  DFFSR \buffer_reg[128]  ( .D(n1316), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[128]) );
  DFFSR \buffer_reg[129]  ( .D(n1315), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[129]) );
  DFFSR \buffer_reg[130]  ( .D(n1314), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[130]) );
  DFFSR \buffer_reg[131]  ( .D(n1313), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[131]) );
  DFFSR \buffer_reg[132]  ( .D(n1312), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[132]) );
  DFFSR \buffer_reg[133]  ( .D(n1311), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[133]) );
  DFFSR \buffer_reg[134]  ( .D(n1310), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[134]) );
  DFFSR \buffer_reg[135]  ( .D(n1309), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[135]) );
  DFFSR \buffer_reg[136]  ( .D(n1308), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[136]) );
  DFFSR \buffer_reg[137]  ( .D(n1307), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[137]) );
  DFFSR \buffer_reg[138]  ( .D(n1306), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[138]) );
  DFFSR \buffer_reg[139]  ( .D(n1305), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[139]) );
  DFFSR \buffer_reg[140]  ( .D(n1304), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[140]) );
  DFFSR \buffer_reg[141]  ( .D(n1303), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[141]) );
  DFFSR \buffer_reg[142]  ( .D(n1302), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[142]) );
  DFFSR \buffer_reg[143]  ( .D(n1301), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[143]) );
  DFFSR \buffer_reg[144]  ( .D(n1300), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[144]) );
  DFFSR \buffer_reg[145]  ( .D(n1299), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[145]) );
  DFFSR \buffer_reg[146]  ( .D(n1298), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[146]) );
  DFFSR \buffer_reg[147]  ( .D(n1297), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[147]) );
  DFFSR \buffer_reg[148]  ( .D(n1296), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[148]) );
  DFFSR \buffer_reg[149]  ( .D(n1295), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[149]) );
  DFFSR \buffer_reg[150]  ( .D(n1294), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[150]) );
  DFFSR \buffer_reg[151]  ( .D(n1293), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[151]) );
  DFFSR \buffer_reg[152]  ( .D(n1292), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[152]) );
  DFFSR \buffer_reg[153]  ( .D(n1291), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[153]) );
  DFFSR \buffer_reg[154]  ( .D(n1290), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[154]) );
  DFFSR \buffer_reg[155]  ( .D(n1289), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[155]) );
  DFFSR \buffer_reg[156]  ( .D(n1288), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[156]) );
  DFFSR \buffer_reg[157]  ( .D(n1287), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[157]) );
  DFFSR \buffer_reg[158]  ( .D(n1286), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[158]) );
  DFFSR \buffer_reg[159]  ( .D(n1285), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[159]) );
  DFFSR \buffer_reg[160]  ( .D(n1284), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[160]) );
  DFFSR \buffer_reg[161]  ( .D(n1283), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[161]) );
  DFFSR \buffer_reg[162]  ( .D(n1282), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[162]) );
  DFFSR \buffer_reg[163]  ( .D(n1281), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[163]) );
  DFFSR \buffer_reg[164]  ( .D(n1280), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[164]) );
  DFFSR \buffer_reg[165]  ( .D(n1279), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[165]) );
  DFFSR \buffer_reg[166]  ( .D(n1278), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[166]) );
  DFFSR \buffer_reg[167]  ( .D(n1277), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[167]) );
  DFFSR \buffer_reg[168]  ( .D(n1276), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[168]) );
  DFFSR \buffer_reg[169]  ( .D(n1275), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[169]) );
  DFFSR \buffer_reg[170]  ( .D(n1274), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[170]) );
  DFFSR \buffer_reg[171]  ( .D(n1273), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[171]) );
  DFFSR \buffer_reg[172]  ( .D(n1272), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[172]) );
  DFFSR \buffer_reg[173]  ( .D(n1271), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[173]) );
  DFFSR \buffer_reg[174]  ( .D(n1270), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[174]) );
  DFFSR \buffer_reg[175]  ( .D(n1269), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[175]) );
  DFFSR \buffer_reg[176]  ( .D(n1268), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[176]) );
  DFFSR \buffer_reg[177]  ( .D(n1267), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[177]) );
  DFFSR \buffer_reg[178]  ( .D(n1266), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[178]) );
  DFFSR \buffer_reg[179]  ( .D(n1265), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[179]) );
  DFFSR \buffer_reg[180]  ( .D(n1264), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[180]) );
  DFFSR \buffer_reg[181]  ( .D(n1263), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[181]) );
  DFFSR \buffer_reg[182]  ( .D(n1262), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[182]) );
  DFFSR \buffer_reg[183]  ( .D(n1261), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[183]) );
  DFFSR \buffer_reg[184]  ( .D(n1260), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[184]) );
  DFFSR \buffer_reg[185]  ( .D(n1259), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[185]) );
  DFFSR \buffer_reg[186]  ( .D(n1258), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[186]) );
  DFFSR \buffer_reg[187]  ( .D(n1257), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[187]) );
  DFFSR \buffer_reg[188]  ( .D(n1256), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[188]) );
  DFFSR \buffer_reg[189]  ( .D(n1255), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[189]) );
  DFFSR \buffer_reg[190]  ( .D(n1254), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[190]) );
  DFFSR \buffer_reg[191]  ( .D(n1253), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[191]) );
  DFFSR \buffer_reg[192]  ( .D(n1252), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[192]) );
  DFFSR \buffer_reg[193]  ( .D(n1251), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[193]) );
  DFFSR \buffer_reg[194]  ( .D(n1250), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[194]) );
  DFFSR \buffer_reg[195]  ( .D(n1249), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[195]) );
  DFFSR \buffer_reg[196]  ( .D(n1248), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[196]) );
  DFFSR \buffer_reg[197]  ( .D(n1247), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[197]) );
  DFFSR \buffer_reg[198]  ( .D(n1246), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[198]) );
  DFFSR \buffer_reg[199]  ( .D(n1245), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[199]) );
  DFFSR \buffer_reg[200]  ( .D(n1244), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[200]) );
  DFFSR \buffer_reg[201]  ( .D(n1243), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[201]) );
  DFFSR \buffer_reg[202]  ( .D(n1242), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[202]) );
  DFFSR \buffer_reg[203]  ( .D(n1241), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[203]) );
  DFFSR \buffer_reg[204]  ( .D(n1240), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[204]) );
  DFFSR \buffer_reg[205]  ( .D(n1239), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[205]) );
  DFFSR \buffer_reg[206]  ( .D(n1238), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[206]) );
  DFFSR \buffer_reg[207]  ( .D(n1237), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[207]) );
  DFFSR \buffer_reg[208]  ( .D(n1236), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[208]) );
  DFFSR \buffer_reg[209]  ( .D(n1235), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[209]) );
  DFFSR \buffer_reg[210]  ( .D(n1234), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[210]) );
  DFFSR \buffer_reg[211]  ( .D(n1233), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[211]) );
  DFFSR \buffer_reg[212]  ( .D(n1232), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[212]) );
  DFFSR \buffer_reg[213]  ( .D(n1231), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[213]) );
  DFFSR \buffer_reg[214]  ( .D(n1230), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[214]) );
  DFFSR \buffer_reg[215]  ( .D(n1229), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[215]) );
  DFFSR \buffer_reg[216]  ( .D(n1228), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[216]) );
  DFFSR \buffer_reg[217]  ( .D(n1227), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[217]) );
  DFFSR \buffer_reg[218]  ( .D(n1226), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[218]) );
  DFFSR \buffer_reg[219]  ( .D(n1225), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[219]) );
  DFFSR \buffer_reg[220]  ( .D(n1224), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[220]) );
  DFFSR \buffer_reg[221]  ( .D(n1223), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[221]) );
  DFFSR \buffer_reg[222]  ( .D(n1222), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[222]) );
  DFFSR \buffer_reg[223]  ( .D(n1221), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[223]) );
  DFFSR \buffer_reg[224]  ( .D(n1220), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[224]) );
  DFFSR \buffer_reg[225]  ( .D(n1219), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[225]) );
  DFFSR \buffer_reg[226]  ( .D(n1218), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[226]) );
  DFFSR \buffer_reg[227]  ( .D(n1217), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[227]) );
  DFFSR \buffer_reg[228]  ( .D(n1216), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[228]) );
  DFFSR \buffer_reg[229]  ( .D(n1215), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[229]) );
  DFFSR \buffer_reg[230]  ( .D(n1214), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[230]) );
  DFFSR \buffer_reg[231]  ( .D(n1213), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[231]) );
  DFFSR \buffer_reg[232]  ( .D(n1212), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[232]) );
  DFFSR \buffer_reg[233]  ( .D(n1211), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[233]) );
  DFFSR \buffer_reg[234]  ( .D(n1210), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[234]) );
  DFFSR \buffer_reg[235]  ( .D(n1209), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[235]) );
  DFFSR \buffer_reg[236]  ( .D(n1208), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[236]) );
  DFFSR \buffer_reg[237]  ( .D(n1207), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[237]) );
  DFFSR \buffer_reg[238]  ( .D(n1206), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[238]) );
  DFFSR \buffer_reg[239]  ( .D(n1205), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[239]) );
  DFFSR \buffer_reg[240]  ( .D(n1204), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[240]) );
  DFFSR \buffer_reg[241]  ( .D(n1203), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[241]) );
  DFFSR \buffer_reg[242]  ( .D(n1202), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[242]) );
  DFFSR \buffer_reg[243]  ( .D(n1201), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[243]) );
  DFFSR \buffer_reg[244]  ( .D(n1200), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[244]) );
  DFFSR \buffer_reg[245]  ( .D(n1199), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[245]) );
  DFFSR \buffer_reg[246]  ( .D(n1198), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[246]) );
  DFFSR \buffer_reg[247]  ( .D(n1197), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[247]) );
  DFFSR \buffer_reg[248]  ( .D(n1196), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[248]) );
  DFFSR \buffer_reg[249]  ( .D(n1195), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[249]) );
  DFFSR \buffer_reg[250]  ( .D(n1194), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[250]) );
  DFFSR \buffer_reg[251]  ( .D(n1193), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[251]) );
  DFFSR \buffer_reg[252]  ( .D(n1192), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[252]) );
  DFFSR \buffer_reg[253]  ( .D(n1191), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[253]) );
  DFFSR \buffer_reg[254]  ( .D(n1190), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[254]) );
  DFFSR \buffer_reg[255]  ( .D(n1189), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[255]) );
  DFFSR \buffer_reg[256]  ( .D(n1188), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[256]) );
  DFFSR \buffer_reg[257]  ( .D(n1187), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[257]) );
  DFFSR \buffer_reg[258]  ( .D(n1186), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[258]) );
  DFFSR \buffer_reg[259]  ( .D(n1185), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[259]) );
  DFFSR \buffer_reg[260]  ( .D(n1184), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[260]) );
  DFFSR \buffer_reg[261]  ( .D(n1183), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[261]) );
  DFFSR \buffer_reg[262]  ( .D(n1182), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[262]) );
  DFFSR \buffer_reg[263]  ( .D(n1181), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[263]) );
  DFFSR \buffer_reg[264]  ( .D(n1180), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[264]) );
  DFFSR \buffer_reg[265]  ( .D(n1179), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[265]) );
  DFFSR \buffer_reg[266]  ( .D(n1178), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[266]) );
  DFFSR \buffer_reg[267]  ( .D(n1177), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[267]) );
  DFFSR \buffer_reg[268]  ( .D(n1176), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[268]) );
  DFFSR \buffer_reg[269]  ( .D(n1175), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[269]) );
  DFFSR \buffer_reg[270]  ( .D(n1174), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[270]) );
  DFFSR \buffer_reg[271]  ( .D(n1173), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[271]) );
  DFFSR \buffer_reg[272]  ( .D(n1172), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[272]) );
  DFFSR \buffer_reg[273]  ( .D(n1171), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[273]) );
  DFFSR \buffer_reg[274]  ( .D(n1170), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[274]) );
  DFFSR \buffer_reg[275]  ( .D(n1169), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[275]) );
  DFFSR \buffer_reg[276]  ( .D(n1168), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[276]) );
  DFFSR \buffer_reg[277]  ( .D(n1167), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[277]) );
  DFFSR \buffer_reg[278]  ( .D(n1166), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[278]) );
  DFFSR \buffer_reg[279]  ( .D(n1165), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[279]) );
  DFFSR \buffer_reg[280]  ( .D(n1164), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[280]) );
  DFFSR \buffer_reg[281]  ( .D(n1163), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[281]) );
  DFFSR \buffer_reg[282]  ( .D(n1162), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[282]) );
  DFFSR \buffer_reg[283]  ( .D(n1161), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[283]) );
  DFFSR \buffer_reg[284]  ( .D(n1160), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[284]) );
  DFFSR \buffer_reg[285]  ( .D(n1159), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[285]) );
  DFFSR \buffer_reg[286]  ( .D(n1158), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[286]) );
  DFFSR \buffer_reg[287]  ( .D(n1157), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[287]) );
  DFFSR \buffer_reg[288]  ( .D(n1156), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[288]) );
  DFFSR \buffer_reg[289]  ( .D(n1155), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[289]) );
  DFFSR \buffer_reg[290]  ( .D(n1154), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[290]) );
  DFFSR \buffer_reg[291]  ( .D(n1153), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[291]) );
  DFFSR \buffer_reg[292]  ( .D(n1152), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[292]) );
  DFFSR \buffer_reg[293]  ( .D(n1151), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[293]) );
  DFFSR \buffer_reg[294]  ( .D(n1150), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[294]) );
  DFFSR \buffer_reg[295]  ( .D(n1149), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[295]) );
  DFFSR \buffer_reg[296]  ( .D(n1148), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[296]) );
  DFFSR \buffer_reg[297]  ( .D(n1147), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[297]) );
  DFFSR \buffer_reg[298]  ( .D(n1146), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[298]) );
  DFFSR \buffer_reg[299]  ( .D(n1145), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[299]) );
  DFFSR \buffer_reg[300]  ( .D(n1144), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[300]) );
  DFFSR \buffer_reg[301]  ( .D(n1143), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[301]) );
  DFFSR \buffer_reg[302]  ( .D(n1142), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[302]) );
  DFFSR \buffer_reg[303]  ( .D(n1141), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[303]) );
  DFFSR \buffer_reg[304]  ( .D(n1140), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[304]) );
  DFFSR \buffer_reg[305]  ( .D(n1139), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[305]) );
  DFFSR \buffer_reg[306]  ( .D(n1138), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[306]) );
  DFFSR \buffer_reg[307]  ( .D(n1137), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[307]) );
  DFFSR \buffer_reg[308]  ( .D(n1136), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[308]) );
  DFFSR \buffer_reg[309]  ( .D(n1135), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[309]) );
  DFFSR \buffer_reg[310]  ( .D(n1134), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[310]) );
  DFFSR \buffer_reg[311]  ( .D(n1133), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[311]) );
  DFFSR \buffer_reg[312]  ( .D(n1132), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[312]) );
  DFFSR \buffer_reg[313]  ( .D(n1131), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[313]) );
  DFFSR \buffer_reg[314]  ( .D(n1130), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[314]) );
  DFFSR \buffer_reg[315]  ( .D(n1129), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[315]) );
  DFFSR \buffer_reg[316]  ( .D(n1128), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[316]) );
  DFFSR \buffer_reg[317]  ( .D(n1127), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[317]) );
  DFFSR \buffer_reg[318]  ( .D(n1126), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[318]) );
  DFFSR \buffer_reg[319]  ( .D(n1125), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[319]) );
  DFFSR \buffer_reg[320]  ( .D(n1124), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[320]) );
  DFFSR \buffer_reg[321]  ( .D(n1123), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[321]) );
  DFFSR \buffer_reg[322]  ( .D(n1122), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[322]) );
  DFFSR \buffer_reg[323]  ( .D(n1121), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[323]) );
  DFFSR \buffer_reg[324]  ( .D(n1120), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[324]) );
  DFFSR \buffer_reg[325]  ( .D(n1119), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[325]) );
  DFFSR \buffer_reg[326]  ( .D(n1118), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[326]) );
  DFFSR \buffer_reg[327]  ( .D(n1117), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[327]) );
  DFFSR \buffer_reg[328]  ( .D(n1116), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[328]) );
  DFFSR \buffer_reg[329]  ( .D(n1115), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[329]) );
  DFFSR \buffer_reg[330]  ( .D(n1114), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[330]) );
  DFFSR \buffer_reg[331]  ( .D(n1113), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[331]) );
  DFFSR \buffer_reg[332]  ( .D(n1112), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[332]) );
  DFFSR \buffer_reg[333]  ( .D(n1111), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[333]) );
  DFFSR \buffer_reg[334]  ( .D(n1110), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[334]) );
  DFFSR \buffer_reg[335]  ( .D(n1109), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[335]) );
  DFFSR \buffer_reg[336]  ( .D(n1108), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[336]) );
  DFFSR \buffer_reg[337]  ( .D(n1107), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[337]) );
  DFFSR \buffer_reg[338]  ( .D(n1106), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[338]) );
  DFFSR \buffer_reg[339]  ( .D(n1105), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[339]) );
  DFFSR \buffer_reg[340]  ( .D(n1104), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[340]) );
  DFFSR \buffer_reg[341]  ( .D(n1103), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[341]) );
  DFFSR \buffer_reg[342]  ( .D(n1102), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[342]) );
  DFFSR \buffer_reg[343]  ( .D(n1101), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[343]) );
  DFFSR \buffer_reg[344]  ( .D(n1100), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[344]) );
  DFFSR \buffer_reg[345]  ( .D(n1099), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[345]) );
  DFFSR \buffer_reg[346]  ( .D(n1098), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[346]) );
  DFFSR \buffer_reg[347]  ( .D(n1097), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[347]) );
  DFFSR \buffer_reg[348]  ( .D(n1096), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[348]) );
  DFFSR \buffer_reg[349]  ( .D(n1095), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[349]) );
  DFFSR \buffer_reg[350]  ( .D(n1094), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[350]) );
  DFFSR \buffer_reg[351]  ( .D(n1093), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[351]) );
  DFFSR \buffer_reg[352]  ( .D(n1092), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[352]) );
  DFFSR \buffer_reg[353]  ( .D(n1091), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[353]) );
  DFFSR \buffer_reg[354]  ( .D(n1090), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[354]) );
  DFFSR \buffer_reg[355]  ( .D(n1089), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[355]) );
  DFFSR \buffer_reg[356]  ( .D(n1088), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[356]) );
  DFFSR \buffer_reg[357]  ( .D(n1087), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[357]) );
  DFFSR \buffer_reg[358]  ( .D(n1086), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        buffer[358]) );
  DFFSR \buffer_reg[359]  ( .D(n1085), .CLK(clk), .R(1'b1), .S(n_rst), .Q(
        serial_out) );
  BUFX2 U363 ( .A(n435), .Y(n400) );
  BUFX2 U364 ( .A(n435), .Y(n401) );
  BUFX2 U365 ( .A(n435), .Y(n402) );
  BUFX2 U366 ( .A(n434), .Y(n403) );
  BUFX2 U367 ( .A(n434), .Y(n404) );
  BUFX2 U368 ( .A(n434), .Y(n405) );
  BUFX2 U369 ( .A(n433), .Y(n406) );
  BUFX2 U370 ( .A(n433), .Y(n407) );
  BUFX2 U371 ( .A(n433), .Y(n408) );
  BUFX2 U372 ( .A(n432), .Y(n409) );
  BUFX2 U373 ( .A(n432), .Y(n410) );
  BUFX2 U374 ( .A(n432), .Y(n411) );
  BUFX2 U375 ( .A(n431), .Y(n412) );
  BUFX2 U376 ( .A(n431), .Y(n413) );
  BUFX2 U377 ( .A(n431), .Y(n414) );
  BUFX2 U378 ( .A(n430), .Y(n415) );
  BUFX2 U379 ( .A(n430), .Y(n416) );
  BUFX2 U380 ( .A(n430), .Y(n417) );
  BUFX2 U381 ( .A(n429), .Y(n418) );
  BUFX2 U382 ( .A(n429), .Y(n419) );
  BUFX2 U383 ( .A(n429), .Y(n420) );
  BUFX2 U384 ( .A(n428), .Y(n421) );
  BUFX2 U385 ( .A(n428), .Y(n422) );
  BUFX2 U386 ( .A(n428), .Y(n423) );
  BUFX2 U387 ( .A(n427), .Y(n424) );
  BUFX2 U388 ( .A(n427), .Y(n425) );
  BUFX2 U389 ( .A(n389), .Y(n387) );
  BUFX2 U390 ( .A(n389), .Y(n386) );
  BUFX2 U391 ( .A(n390), .Y(n385) );
  BUFX2 U392 ( .A(n390), .Y(n384) );
  BUFX2 U393 ( .A(n390), .Y(n383) );
  BUFX2 U394 ( .A(n391), .Y(n382) );
  BUFX2 U395 ( .A(n391), .Y(n381) );
  BUFX2 U396 ( .A(n391), .Y(n380) );
  BUFX2 U397 ( .A(n392), .Y(n379) );
  BUFX2 U398 ( .A(n392), .Y(n378) );
  BUFX2 U399 ( .A(n392), .Y(n377) );
  BUFX2 U400 ( .A(n393), .Y(n376) );
  BUFX2 U401 ( .A(n393), .Y(n375) );
  BUFX2 U402 ( .A(n393), .Y(n374) );
  BUFX2 U403 ( .A(n394), .Y(n373) );
  BUFX2 U404 ( .A(n394), .Y(n372) );
  BUFX2 U405 ( .A(n394), .Y(n371) );
  BUFX2 U406 ( .A(n395), .Y(n370) );
  BUFX2 U407 ( .A(n395), .Y(n369) );
  BUFX2 U408 ( .A(n395), .Y(n368) );
  BUFX2 U409 ( .A(n396), .Y(n367) );
  BUFX2 U410 ( .A(n396), .Y(n366) );
  BUFX2 U411 ( .A(n396), .Y(n365) );
  BUFX2 U412 ( .A(n397), .Y(n364) );
  BUFX2 U413 ( .A(n397), .Y(n363) );
  BUFX2 U414 ( .A(n397), .Y(n362) );
  BUFX2 U415 ( .A(n389), .Y(n388) );
  BUFX2 U416 ( .A(n427), .Y(n426) );
  BUFX2 U417 ( .A(n436), .Y(n399) );
  BUFX2 U418 ( .A(n478), .Y(n436) );
  BUFX2 U419 ( .A(n398), .Y(n361) );
  BUFX2 U420 ( .A(n476), .Y(n398) );
  BUFX2 U421 ( .A(n478), .Y(n435) );
  BUFX2 U422 ( .A(n478), .Y(n434) );
  BUFX2 U423 ( .A(n478), .Y(n433) );
  BUFX2 U424 ( .A(n478), .Y(n432) );
  BUFX2 U425 ( .A(n478), .Y(n431) );
  BUFX2 U426 ( .A(n478), .Y(n430) );
  BUFX2 U427 ( .A(n478), .Y(n429) );
  BUFX2 U428 ( .A(n478), .Y(n428) );
  BUFX2 U429 ( .A(n478), .Y(n427) );
  BUFX2 U430 ( .A(n476), .Y(n389) );
  BUFX2 U431 ( .A(n476), .Y(n390) );
  BUFX2 U432 ( .A(n476), .Y(n391) );
  BUFX2 U433 ( .A(n476), .Y(n392) );
  BUFX2 U434 ( .A(n476), .Y(n393) );
  BUFX2 U435 ( .A(n476), .Y(n394) );
  BUFX2 U436 ( .A(n476), .Y(n395) );
  BUFX2 U437 ( .A(n476), .Y(n396) );
  BUFX2 U438 ( .A(n476), .Y(n397) );
  BUFX2 U439 ( .A(n469), .Y(n451) );
  BUFX2 U440 ( .A(n469), .Y(n452) );
  BUFX2 U441 ( .A(n468), .Y(n453) );
  BUFX2 U442 ( .A(n468), .Y(n454) );
  BUFX2 U443 ( .A(n468), .Y(n455) );
  BUFX2 U444 ( .A(n467), .Y(n456) );
  BUFX2 U445 ( .A(n467), .Y(n457) );
  BUFX2 U446 ( .A(n467), .Y(n458) );
  BUFX2 U447 ( .A(n466), .Y(n459) );
  BUFX2 U448 ( .A(n466), .Y(n460) );
  BUFX2 U449 ( .A(n466), .Y(n461) );
  BUFX2 U450 ( .A(n465), .Y(n462) );
  BUFX2 U451 ( .A(n465), .Y(n463) );
  BUFX2 U452 ( .A(n473), .Y(n438) );
  BUFX2 U453 ( .A(n473), .Y(n439) );
  BUFX2 U454 ( .A(n473), .Y(n440) );
  BUFX2 U455 ( .A(n472), .Y(n441) );
  BUFX2 U456 ( .A(n472), .Y(n442) );
  BUFX2 U457 ( .A(n472), .Y(n443) );
  BUFX2 U458 ( .A(n471), .Y(n444) );
  BUFX2 U459 ( .A(n471), .Y(n445) );
  BUFX2 U460 ( .A(n471), .Y(n446) );
  BUFX2 U461 ( .A(n470), .Y(n447) );
  BUFX2 U462 ( .A(n470), .Y(n448) );
  BUFX2 U463 ( .A(n470), .Y(n449) );
  BUFX2 U464 ( .A(n469), .Y(n450) );
  BUFX2 U465 ( .A(n465), .Y(n464) );
  BUFX2 U466 ( .A(n474), .Y(n437) );
  BUFX2 U467 ( .A(n479), .Y(n474) );
  BUFX2 U468 ( .A(n479), .Y(n468) );
  BUFX2 U469 ( .A(n479), .Y(n467) );
  BUFX2 U470 ( .A(n479), .Y(n466) );
  BUFX2 U471 ( .A(n479), .Y(n465) );
  BUFX2 U472 ( .A(n479), .Y(n473) );
  BUFX2 U473 ( .A(n479), .Y(n472) );
  BUFX2 U474 ( .A(n479), .Y(n471) );
  BUFX2 U475 ( .A(n479), .Y(n470) );
  BUFX2 U476 ( .A(n479), .Y(n469) );
  OAI21X1 U477 ( .A(n475), .B(n361), .C(n477), .Y(n1444) );
  AOI21X1 U478 ( .A(n426), .B(buffer[0]), .C(n464), .Y(n477) );
  INVX1 U479 ( .A(parallel_in[0]), .Y(n475) );
  OAI21X1 U480 ( .A(n361), .B(n480), .C(n481), .Y(n1443) );
  AOI22X1 U481 ( .A(buffer[1]), .B(n426), .C(n464), .D(buffer[0]), .Y(n481) );
  INVX1 U482 ( .A(parallel_in[1]), .Y(n480) );
  OAI21X1 U483 ( .A(n361), .B(n482), .C(n483), .Y(n1442) );
  AOI22X1 U484 ( .A(buffer[2]), .B(n426), .C(n464), .D(buffer[1]), .Y(n483) );
  INVX1 U485 ( .A(parallel_in[2]), .Y(n482) );
  OAI21X1 U486 ( .A(n361), .B(n484), .C(n485), .Y(n1441) );
  AOI22X1 U487 ( .A(buffer[3]), .B(n426), .C(buffer[2]), .D(n437), .Y(n485) );
  INVX1 U488 ( .A(parallel_in[3]), .Y(n484) );
  OAI21X1 U489 ( .A(n361), .B(n486), .C(n487), .Y(n1440) );
  AOI22X1 U490 ( .A(buffer[4]), .B(n426), .C(buffer[3]), .D(n450), .Y(n487) );
  INVX1 U491 ( .A(parallel_in[4]), .Y(n486) );
  OAI21X1 U492 ( .A(n361), .B(n488), .C(n489), .Y(n1439) );
  AOI22X1 U493 ( .A(buffer[5]), .B(n426), .C(buffer[4]), .D(n450), .Y(n489) );
  INVX1 U494 ( .A(parallel_in[5]), .Y(n488) );
  OAI21X1 U495 ( .A(n361), .B(n490), .C(n491), .Y(n1438) );
  AOI22X1 U496 ( .A(buffer[6]), .B(n426), .C(buffer[5]), .D(n450), .Y(n491) );
  INVX1 U497 ( .A(parallel_in[6]), .Y(n490) );
  OAI21X1 U498 ( .A(n361), .B(n492), .C(n493), .Y(n1437) );
  AOI22X1 U499 ( .A(buffer[7]), .B(n426), .C(buffer[6]), .D(n450), .Y(n493) );
  INVX1 U500 ( .A(parallel_in[7]), .Y(n492) );
  OAI21X1 U501 ( .A(n361), .B(n494), .C(n495), .Y(n1436) );
  AOI22X1 U502 ( .A(buffer[8]), .B(n426), .C(buffer[7]), .D(n450), .Y(n495) );
  INVX1 U503 ( .A(parallel_in[8]), .Y(n494) );
  OAI21X1 U504 ( .A(n361), .B(n496), .C(n497), .Y(n1435) );
  AOI22X1 U505 ( .A(buffer[9]), .B(n425), .C(buffer[8]), .D(n450), .Y(n497) );
  INVX1 U506 ( .A(parallel_in[9]), .Y(n496) );
  OAI21X1 U507 ( .A(n361), .B(n498), .C(n499), .Y(n1434) );
  AOI22X1 U508 ( .A(buffer[10]), .B(n425), .C(buffer[9]), .D(n450), .Y(n499)
         );
  INVX1 U509 ( .A(parallel_in[10]), .Y(n498) );
  OAI21X1 U510 ( .A(n361), .B(n500), .C(n501), .Y(n1433) );
  AOI22X1 U511 ( .A(buffer[11]), .B(n425), .C(buffer[10]), .D(n450), .Y(n501)
         );
  INVX1 U512 ( .A(parallel_in[11]), .Y(n500) );
  OAI21X1 U513 ( .A(n361), .B(n502), .C(n503), .Y(n1432) );
  AOI22X1 U514 ( .A(buffer[12]), .B(n425), .C(buffer[11]), .D(n450), .Y(n503)
         );
  INVX1 U515 ( .A(parallel_in[12]), .Y(n502) );
  OAI21X1 U516 ( .A(n362), .B(n504), .C(n505), .Y(n1431) );
  AOI22X1 U517 ( .A(buffer[13]), .B(n425), .C(buffer[12]), .D(n449), .Y(n505)
         );
  INVX1 U518 ( .A(parallel_in[13]), .Y(n504) );
  OAI21X1 U519 ( .A(n362), .B(n506), .C(n507), .Y(n1430) );
  AOI22X1 U520 ( .A(buffer[14]), .B(n425), .C(buffer[13]), .D(n449), .Y(n507)
         );
  INVX1 U521 ( .A(parallel_in[14]), .Y(n506) );
  OAI21X1 U522 ( .A(n362), .B(n508), .C(n509), .Y(n1429) );
  AOI22X1 U523 ( .A(buffer[15]), .B(n425), .C(buffer[14]), .D(n449), .Y(n509)
         );
  INVX1 U524 ( .A(parallel_in[15]), .Y(n508) );
  OAI21X1 U525 ( .A(n362), .B(n510), .C(n511), .Y(n1428) );
  AOI22X1 U526 ( .A(buffer[16]), .B(n425), .C(buffer[15]), .D(n449), .Y(n511)
         );
  INVX1 U527 ( .A(parallel_in[16]), .Y(n510) );
  OAI21X1 U528 ( .A(n362), .B(n512), .C(n513), .Y(n1427) );
  AOI22X1 U529 ( .A(buffer[17]), .B(n425), .C(buffer[16]), .D(n449), .Y(n513)
         );
  INVX1 U530 ( .A(parallel_in[17]), .Y(n512) );
  OAI21X1 U531 ( .A(n362), .B(n514), .C(n515), .Y(n1426) );
  AOI22X1 U532 ( .A(buffer[18]), .B(n425), .C(buffer[17]), .D(n449), .Y(n515)
         );
  INVX1 U533 ( .A(parallel_in[18]), .Y(n514) );
  OAI21X1 U534 ( .A(n362), .B(n516), .C(n517), .Y(n1425) );
  AOI22X1 U535 ( .A(buffer[19]), .B(n425), .C(buffer[18]), .D(n449), .Y(n517)
         );
  INVX1 U536 ( .A(parallel_in[19]), .Y(n516) );
  OAI21X1 U537 ( .A(n362), .B(n518), .C(n519), .Y(n1424) );
  AOI22X1 U538 ( .A(buffer[20]), .B(n425), .C(buffer[19]), .D(n449), .Y(n519)
         );
  INVX1 U539 ( .A(parallel_in[20]), .Y(n518) );
  OAI21X1 U540 ( .A(n362), .B(n520), .C(n521), .Y(n1423) );
  AOI22X1 U541 ( .A(buffer[21]), .B(n425), .C(buffer[20]), .D(n449), .Y(n521)
         );
  INVX1 U542 ( .A(parallel_in[21]), .Y(n520) );
  OAI21X1 U543 ( .A(n362), .B(n522), .C(n523), .Y(n1422) );
  AOI22X1 U544 ( .A(buffer[22]), .B(n424), .C(buffer[21]), .D(n449), .Y(n523)
         );
  INVX1 U545 ( .A(parallel_in[22]), .Y(n522) );
  OAI21X1 U546 ( .A(n362), .B(n524), .C(n525), .Y(n1421) );
  AOI22X1 U547 ( .A(buffer[23]), .B(n424), .C(buffer[22]), .D(n449), .Y(n525)
         );
  INVX1 U548 ( .A(parallel_in[23]), .Y(n524) );
  OAI21X1 U549 ( .A(n362), .B(n526), .C(n527), .Y(n1420) );
  AOI22X1 U550 ( .A(buffer[24]), .B(n424), .C(buffer[23]), .D(n449), .Y(n527)
         );
  INVX1 U551 ( .A(parallel_in[24]), .Y(n526) );
  OAI21X1 U552 ( .A(n362), .B(n528), .C(n529), .Y(n1419) );
  AOI22X1 U553 ( .A(buffer[25]), .B(n424), .C(buffer[24]), .D(n449), .Y(n529)
         );
  INVX1 U554 ( .A(parallel_in[25]), .Y(n528) );
  OAI21X1 U555 ( .A(n363), .B(n530), .C(n531), .Y(n1418) );
  AOI22X1 U556 ( .A(buffer[26]), .B(n424), .C(buffer[25]), .D(n448), .Y(n531)
         );
  INVX1 U557 ( .A(parallel_in[26]), .Y(n530) );
  OAI21X1 U558 ( .A(n363), .B(n532), .C(n533), .Y(n1417) );
  AOI22X1 U559 ( .A(buffer[27]), .B(n424), .C(buffer[26]), .D(n448), .Y(n533)
         );
  INVX1 U560 ( .A(parallel_in[27]), .Y(n532) );
  OAI21X1 U561 ( .A(n363), .B(n534), .C(n535), .Y(n1416) );
  AOI22X1 U562 ( .A(buffer[28]), .B(n424), .C(buffer[27]), .D(n448), .Y(n535)
         );
  INVX1 U563 ( .A(parallel_in[28]), .Y(n534) );
  OAI21X1 U564 ( .A(n363), .B(n536), .C(n537), .Y(n1415) );
  AOI22X1 U565 ( .A(buffer[29]), .B(n424), .C(buffer[28]), .D(n448), .Y(n537)
         );
  INVX1 U566 ( .A(parallel_in[29]), .Y(n536) );
  OAI21X1 U567 ( .A(n363), .B(n538), .C(n539), .Y(n1414) );
  AOI22X1 U568 ( .A(buffer[30]), .B(n424), .C(buffer[29]), .D(n448), .Y(n539)
         );
  INVX1 U569 ( .A(parallel_in[30]), .Y(n538) );
  OAI21X1 U570 ( .A(n363), .B(n540), .C(n541), .Y(n1413) );
  AOI22X1 U571 ( .A(buffer[31]), .B(n424), .C(buffer[30]), .D(n448), .Y(n541)
         );
  INVX1 U572 ( .A(parallel_in[31]), .Y(n540) );
  OAI21X1 U573 ( .A(n363), .B(n542), .C(n543), .Y(n1412) );
  AOI22X1 U574 ( .A(buffer[32]), .B(n424), .C(buffer[31]), .D(n448), .Y(n543)
         );
  INVX1 U575 ( .A(parallel_in[32]), .Y(n542) );
  OAI21X1 U576 ( .A(n363), .B(n544), .C(n545), .Y(n1411) );
  AOI22X1 U577 ( .A(buffer[33]), .B(n424), .C(buffer[32]), .D(n448), .Y(n545)
         );
  INVX1 U578 ( .A(parallel_in[33]), .Y(n544) );
  OAI21X1 U579 ( .A(n363), .B(n546), .C(n547), .Y(n1410) );
  AOI22X1 U580 ( .A(buffer[34]), .B(n424), .C(buffer[33]), .D(n448), .Y(n547)
         );
  INVX1 U581 ( .A(parallel_in[34]), .Y(n546) );
  OAI21X1 U582 ( .A(n363), .B(n548), .C(n549), .Y(n1409) );
  AOI22X1 U583 ( .A(buffer[35]), .B(n423), .C(buffer[34]), .D(n448), .Y(n549)
         );
  INVX1 U584 ( .A(parallel_in[35]), .Y(n548) );
  OAI21X1 U585 ( .A(n363), .B(n550), .C(n551), .Y(n1408) );
  AOI22X1 U586 ( .A(buffer[36]), .B(n423), .C(buffer[35]), .D(n448), .Y(n551)
         );
  INVX1 U587 ( .A(parallel_in[36]), .Y(n550) );
  OAI21X1 U588 ( .A(n363), .B(n552), .C(n553), .Y(n1407) );
  AOI22X1 U589 ( .A(buffer[37]), .B(n423), .C(buffer[36]), .D(n448), .Y(n553)
         );
  INVX1 U590 ( .A(parallel_in[37]), .Y(n552) );
  OAI21X1 U591 ( .A(n363), .B(n554), .C(n555), .Y(n1406) );
  AOI22X1 U592 ( .A(buffer[38]), .B(n423), .C(buffer[37]), .D(n448), .Y(n555)
         );
  INVX1 U593 ( .A(parallel_in[38]), .Y(n554) );
  OAI21X1 U594 ( .A(n364), .B(n556), .C(n557), .Y(n1405) );
  AOI22X1 U595 ( .A(buffer[39]), .B(n423), .C(buffer[38]), .D(n447), .Y(n557)
         );
  INVX1 U596 ( .A(parallel_in[39]), .Y(n556) );
  OAI21X1 U597 ( .A(n364), .B(n558), .C(n559), .Y(n1404) );
  AOI22X1 U598 ( .A(buffer[40]), .B(n423), .C(buffer[39]), .D(n447), .Y(n559)
         );
  INVX1 U599 ( .A(parallel_in[40]), .Y(n558) );
  OAI21X1 U600 ( .A(n364), .B(n560), .C(n561), .Y(n1403) );
  AOI22X1 U601 ( .A(buffer[41]), .B(n423), .C(buffer[40]), .D(n447), .Y(n561)
         );
  INVX1 U602 ( .A(parallel_in[41]), .Y(n560) );
  OAI21X1 U603 ( .A(n364), .B(n562), .C(n563), .Y(n1402) );
  AOI22X1 U604 ( .A(buffer[42]), .B(n423), .C(buffer[41]), .D(n447), .Y(n563)
         );
  INVX1 U605 ( .A(parallel_in[42]), .Y(n562) );
  OAI21X1 U606 ( .A(n364), .B(n564), .C(n565), .Y(n1401) );
  AOI22X1 U607 ( .A(buffer[43]), .B(n423), .C(buffer[42]), .D(n447), .Y(n565)
         );
  INVX1 U608 ( .A(parallel_in[43]), .Y(n564) );
  OAI21X1 U609 ( .A(n364), .B(n566), .C(n567), .Y(n1400) );
  AOI22X1 U610 ( .A(buffer[44]), .B(n423), .C(buffer[43]), .D(n447), .Y(n567)
         );
  INVX1 U611 ( .A(parallel_in[44]), .Y(n566) );
  OAI21X1 U612 ( .A(n364), .B(n568), .C(n569), .Y(n1399) );
  AOI22X1 U613 ( .A(buffer[45]), .B(n423), .C(buffer[44]), .D(n447), .Y(n569)
         );
  INVX1 U614 ( .A(parallel_in[45]), .Y(n568) );
  OAI21X1 U615 ( .A(n364), .B(n570), .C(n571), .Y(n1398) );
  AOI22X1 U616 ( .A(buffer[46]), .B(n423), .C(buffer[45]), .D(n447), .Y(n571)
         );
  INVX1 U617 ( .A(parallel_in[46]), .Y(n570) );
  OAI21X1 U618 ( .A(n364), .B(n572), .C(n573), .Y(n1397) );
  AOI22X1 U619 ( .A(buffer[47]), .B(n423), .C(buffer[46]), .D(n447), .Y(n573)
         );
  INVX1 U620 ( .A(parallel_in[47]), .Y(n572) );
  OAI21X1 U621 ( .A(n364), .B(n574), .C(n575), .Y(n1396) );
  AOI22X1 U622 ( .A(buffer[48]), .B(n422), .C(buffer[47]), .D(n447), .Y(n575)
         );
  INVX1 U623 ( .A(parallel_in[48]), .Y(n574) );
  OAI21X1 U624 ( .A(n364), .B(n576), .C(n577), .Y(n1395) );
  AOI22X1 U625 ( .A(buffer[49]), .B(n422), .C(buffer[48]), .D(n447), .Y(n577)
         );
  INVX1 U626 ( .A(parallel_in[49]), .Y(n576) );
  OAI21X1 U627 ( .A(n364), .B(n578), .C(n579), .Y(n1394) );
  AOI22X1 U628 ( .A(buffer[50]), .B(n422), .C(buffer[49]), .D(n447), .Y(n579)
         );
  INVX1 U629 ( .A(parallel_in[50]), .Y(n578) );
  OAI21X1 U630 ( .A(n364), .B(n580), .C(n581), .Y(n1393) );
  AOI22X1 U631 ( .A(buffer[51]), .B(n422), .C(buffer[50]), .D(n447), .Y(n581)
         );
  INVX1 U632 ( .A(parallel_in[51]), .Y(n580) );
  OAI21X1 U633 ( .A(n365), .B(n582), .C(n583), .Y(n1392) );
  AOI22X1 U634 ( .A(buffer[52]), .B(n422), .C(buffer[51]), .D(n446), .Y(n583)
         );
  INVX1 U635 ( .A(parallel_in[52]), .Y(n582) );
  OAI21X1 U636 ( .A(n365), .B(n584), .C(n585), .Y(n1391) );
  AOI22X1 U637 ( .A(buffer[53]), .B(n422), .C(buffer[52]), .D(n446), .Y(n585)
         );
  INVX1 U638 ( .A(parallel_in[53]), .Y(n584) );
  OAI21X1 U639 ( .A(n365), .B(n586), .C(n587), .Y(n1390) );
  AOI22X1 U640 ( .A(buffer[54]), .B(n422), .C(buffer[53]), .D(n446), .Y(n587)
         );
  INVX1 U641 ( .A(parallel_in[54]), .Y(n586) );
  OAI21X1 U642 ( .A(n365), .B(n588), .C(n589), .Y(n1389) );
  AOI22X1 U643 ( .A(buffer[55]), .B(n422), .C(buffer[54]), .D(n446), .Y(n589)
         );
  INVX1 U644 ( .A(parallel_in[55]), .Y(n588) );
  OAI21X1 U645 ( .A(n365), .B(n590), .C(n591), .Y(n1388) );
  AOI22X1 U646 ( .A(buffer[56]), .B(n422), .C(buffer[55]), .D(n446), .Y(n591)
         );
  INVX1 U647 ( .A(parallel_in[56]), .Y(n590) );
  OAI21X1 U648 ( .A(n365), .B(n592), .C(n593), .Y(n1387) );
  AOI22X1 U649 ( .A(buffer[57]), .B(n422), .C(buffer[56]), .D(n446), .Y(n593)
         );
  INVX1 U650 ( .A(parallel_in[57]), .Y(n592) );
  OAI21X1 U651 ( .A(n365), .B(n594), .C(n595), .Y(n1386) );
  AOI22X1 U652 ( .A(buffer[58]), .B(n422), .C(buffer[57]), .D(n446), .Y(n595)
         );
  INVX1 U653 ( .A(parallel_in[58]), .Y(n594) );
  OAI21X1 U654 ( .A(n365), .B(n596), .C(n597), .Y(n1385) );
  AOI22X1 U655 ( .A(buffer[59]), .B(n422), .C(buffer[58]), .D(n446), .Y(n597)
         );
  INVX1 U656 ( .A(parallel_in[59]), .Y(n596) );
  OAI21X1 U657 ( .A(n365), .B(n598), .C(n599), .Y(n1384) );
  AOI22X1 U658 ( .A(buffer[60]), .B(n422), .C(buffer[59]), .D(n446), .Y(n599)
         );
  INVX1 U659 ( .A(parallel_in[60]), .Y(n598) );
  OAI21X1 U660 ( .A(n365), .B(n600), .C(n601), .Y(n1383) );
  AOI22X1 U661 ( .A(buffer[61]), .B(n421), .C(buffer[60]), .D(n446), .Y(n601)
         );
  INVX1 U662 ( .A(parallel_in[61]), .Y(n600) );
  OAI21X1 U663 ( .A(n365), .B(n602), .C(n603), .Y(n1382) );
  AOI22X1 U664 ( .A(buffer[62]), .B(n421), .C(buffer[61]), .D(n446), .Y(n603)
         );
  INVX1 U665 ( .A(parallel_in[62]), .Y(n602) );
  OAI21X1 U666 ( .A(n365), .B(n604), .C(n605), .Y(n1381) );
  AOI22X1 U667 ( .A(buffer[63]), .B(n421), .C(buffer[62]), .D(n446), .Y(n605)
         );
  INVX1 U668 ( .A(parallel_in[63]), .Y(n604) );
  OAI21X1 U669 ( .A(n365), .B(n606), .C(n607), .Y(n1380) );
  AOI22X1 U670 ( .A(buffer[64]), .B(n421), .C(buffer[63]), .D(n446), .Y(n607)
         );
  INVX1 U671 ( .A(parallel_in[64]), .Y(n606) );
  OAI21X1 U672 ( .A(n366), .B(n608), .C(n609), .Y(n1379) );
  AOI22X1 U673 ( .A(buffer[65]), .B(n421), .C(buffer[64]), .D(n445), .Y(n609)
         );
  INVX1 U674 ( .A(parallel_in[65]), .Y(n608) );
  OAI21X1 U675 ( .A(n366), .B(n610), .C(n611), .Y(n1378) );
  AOI22X1 U676 ( .A(buffer[66]), .B(n421), .C(buffer[65]), .D(n445), .Y(n611)
         );
  INVX1 U677 ( .A(parallel_in[66]), .Y(n610) );
  OAI21X1 U678 ( .A(n366), .B(n612), .C(n613), .Y(n1377) );
  AOI22X1 U679 ( .A(buffer[67]), .B(n421), .C(buffer[66]), .D(n445), .Y(n613)
         );
  INVX1 U680 ( .A(parallel_in[67]), .Y(n612) );
  OAI21X1 U681 ( .A(n366), .B(n614), .C(n615), .Y(n1376) );
  AOI22X1 U682 ( .A(buffer[68]), .B(n421), .C(buffer[67]), .D(n445), .Y(n615)
         );
  INVX1 U683 ( .A(parallel_in[68]), .Y(n614) );
  OAI21X1 U684 ( .A(n366), .B(n616), .C(n617), .Y(n1375) );
  AOI22X1 U685 ( .A(buffer[69]), .B(n421), .C(buffer[68]), .D(n445), .Y(n617)
         );
  INVX1 U686 ( .A(parallel_in[69]), .Y(n616) );
  OAI21X1 U687 ( .A(n366), .B(n618), .C(n619), .Y(n1374) );
  AOI22X1 U688 ( .A(buffer[70]), .B(n421), .C(buffer[69]), .D(n445), .Y(n619)
         );
  INVX1 U689 ( .A(parallel_in[70]), .Y(n618) );
  OAI21X1 U690 ( .A(n366), .B(n620), .C(n621), .Y(n1373) );
  AOI22X1 U691 ( .A(buffer[71]), .B(n421), .C(buffer[70]), .D(n445), .Y(n621)
         );
  INVX1 U692 ( .A(parallel_in[71]), .Y(n620) );
  OAI21X1 U693 ( .A(n366), .B(n622), .C(n623), .Y(n1372) );
  AOI22X1 U694 ( .A(buffer[72]), .B(n421), .C(buffer[71]), .D(n445), .Y(n623)
         );
  INVX1 U695 ( .A(parallel_in[72]), .Y(n622) );
  OAI21X1 U696 ( .A(n366), .B(n624), .C(n625), .Y(n1371) );
  AOI22X1 U697 ( .A(buffer[73]), .B(n421), .C(buffer[72]), .D(n445), .Y(n625)
         );
  INVX1 U698 ( .A(parallel_in[73]), .Y(n624) );
  OAI21X1 U699 ( .A(n366), .B(n626), .C(n627), .Y(n1370) );
  AOI22X1 U700 ( .A(buffer[74]), .B(n420), .C(buffer[73]), .D(n445), .Y(n627)
         );
  INVX1 U701 ( .A(parallel_in[74]), .Y(n626) );
  OAI21X1 U702 ( .A(n366), .B(n628), .C(n629), .Y(n1369) );
  AOI22X1 U703 ( .A(buffer[75]), .B(n420), .C(buffer[74]), .D(n445), .Y(n629)
         );
  INVX1 U704 ( .A(parallel_in[75]), .Y(n628) );
  OAI21X1 U705 ( .A(n366), .B(n630), .C(n631), .Y(n1368) );
  AOI22X1 U706 ( .A(buffer[76]), .B(n420), .C(buffer[75]), .D(n445), .Y(n631)
         );
  INVX1 U707 ( .A(parallel_in[76]), .Y(n630) );
  OAI21X1 U708 ( .A(n366), .B(n632), .C(n633), .Y(n1367) );
  AOI22X1 U709 ( .A(buffer[77]), .B(n420), .C(buffer[76]), .D(n445), .Y(n633)
         );
  INVX1 U710 ( .A(parallel_in[77]), .Y(n632) );
  OAI21X1 U711 ( .A(n367), .B(n634), .C(n635), .Y(n1366) );
  AOI22X1 U712 ( .A(buffer[78]), .B(n420), .C(buffer[77]), .D(n444), .Y(n635)
         );
  INVX1 U713 ( .A(parallel_in[78]), .Y(n634) );
  OAI21X1 U714 ( .A(n367), .B(n636), .C(n637), .Y(n1365) );
  AOI22X1 U715 ( .A(buffer[79]), .B(n420), .C(buffer[78]), .D(n444), .Y(n637)
         );
  INVX1 U716 ( .A(parallel_in[79]), .Y(n636) );
  OAI21X1 U717 ( .A(n367), .B(n638), .C(n639), .Y(n1364) );
  AOI22X1 U718 ( .A(buffer[80]), .B(n420), .C(buffer[79]), .D(n444), .Y(n639)
         );
  INVX1 U719 ( .A(parallel_in[80]), .Y(n638) );
  OAI21X1 U720 ( .A(n367), .B(n640), .C(n641), .Y(n1363) );
  AOI22X1 U721 ( .A(buffer[81]), .B(n420), .C(buffer[80]), .D(n444), .Y(n641)
         );
  INVX1 U722 ( .A(parallel_in[81]), .Y(n640) );
  OAI21X1 U723 ( .A(n367), .B(n642), .C(n643), .Y(n1362) );
  AOI22X1 U724 ( .A(buffer[82]), .B(n420), .C(buffer[81]), .D(n444), .Y(n643)
         );
  INVX1 U725 ( .A(parallel_in[82]), .Y(n642) );
  OAI21X1 U726 ( .A(n367), .B(n644), .C(n645), .Y(n1361) );
  AOI22X1 U727 ( .A(buffer[83]), .B(n420), .C(buffer[82]), .D(n444), .Y(n645)
         );
  INVX1 U728 ( .A(parallel_in[83]), .Y(n644) );
  OAI21X1 U729 ( .A(n367), .B(n646), .C(n647), .Y(n1360) );
  AOI22X1 U730 ( .A(buffer[84]), .B(n420), .C(buffer[83]), .D(n444), .Y(n647)
         );
  INVX1 U731 ( .A(parallel_in[84]), .Y(n646) );
  OAI21X1 U732 ( .A(n367), .B(n648), .C(n649), .Y(n1359) );
  AOI22X1 U733 ( .A(buffer[85]), .B(n420), .C(buffer[84]), .D(n444), .Y(n649)
         );
  INVX1 U734 ( .A(parallel_in[85]), .Y(n648) );
  OAI21X1 U735 ( .A(n367), .B(n650), .C(n651), .Y(n1358) );
  AOI22X1 U736 ( .A(buffer[86]), .B(n420), .C(buffer[85]), .D(n444), .Y(n651)
         );
  INVX1 U737 ( .A(parallel_in[86]), .Y(n650) );
  OAI21X1 U738 ( .A(n367), .B(n652), .C(n653), .Y(n1357) );
  AOI22X1 U739 ( .A(buffer[87]), .B(n419), .C(buffer[86]), .D(n444), .Y(n653)
         );
  INVX1 U740 ( .A(parallel_in[87]), .Y(n652) );
  OAI21X1 U741 ( .A(n367), .B(n654), .C(n655), .Y(n1356) );
  AOI22X1 U742 ( .A(buffer[88]), .B(n419), .C(buffer[87]), .D(n444), .Y(n655)
         );
  INVX1 U743 ( .A(parallel_in[88]), .Y(n654) );
  OAI21X1 U744 ( .A(n367), .B(n656), .C(n657), .Y(n1355) );
  AOI22X1 U745 ( .A(buffer[89]), .B(n419), .C(buffer[88]), .D(n444), .Y(n657)
         );
  INVX1 U746 ( .A(parallel_in[89]), .Y(n656) );
  OAI21X1 U747 ( .A(n367), .B(n658), .C(n659), .Y(n1354) );
  AOI22X1 U748 ( .A(buffer[90]), .B(n419), .C(buffer[89]), .D(n450), .Y(n659)
         );
  INVX1 U749 ( .A(parallel_in[90]), .Y(n658) );
  OAI21X1 U750 ( .A(n368), .B(n660), .C(n661), .Y(n1353) );
  AOI22X1 U751 ( .A(buffer[91]), .B(n419), .C(buffer[90]), .D(n444), .Y(n661)
         );
  INVX1 U752 ( .A(parallel_in[91]), .Y(n660) );
  OAI21X1 U753 ( .A(n368), .B(n662), .C(n663), .Y(n1352) );
  AOI22X1 U754 ( .A(buffer[92]), .B(n419), .C(buffer[91]), .D(n443), .Y(n663)
         );
  INVX1 U755 ( .A(parallel_in[92]), .Y(n662) );
  OAI21X1 U756 ( .A(n368), .B(n664), .C(n665), .Y(n1351) );
  AOI22X1 U757 ( .A(buffer[93]), .B(n419), .C(buffer[92]), .D(n443), .Y(n665)
         );
  INVX1 U758 ( .A(parallel_in[93]), .Y(n664) );
  OAI21X1 U759 ( .A(n368), .B(n666), .C(n667), .Y(n1350) );
  AOI22X1 U760 ( .A(buffer[94]), .B(n419), .C(buffer[93]), .D(n443), .Y(n667)
         );
  INVX1 U761 ( .A(parallel_in[94]), .Y(n666) );
  OAI21X1 U762 ( .A(n368), .B(n668), .C(n669), .Y(n1349) );
  AOI22X1 U763 ( .A(buffer[95]), .B(n419), .C(buffer[94]), .D(n443), .Y(n669)
         );
  INVX1 U764 ( .A(parallel_in[95]), .Y(n668) );
  OAI21X1 U765 ( .A(n368), .B(n670), .C(n671), .Y(n1348) );
  AOI22X1 U766 ( .A(buffer[96]), .B(n419), .C(buffer[95]), .D(n443), .Y(n671)
         );
  INVX1 U767 ( .A(parallel_in[96]), .Y(n670) );
  OAI21X1 U768 ( .A(n368), .B(n672), .C(n673), .Y(n1347) );
  AOI22X1 U769 ( .A(buffer[97]), .B(n419), .C(buffer[96]), .D(n443), .Y(n673)
         );
  INVX1 U770 ( .A(parallel_in[97]), .Y(n672) );
  OAI21X1 U771 ( .A(n368), .B(n674), .C(n675), .Y(n1346) );
  AOI22X1 U772 ( .A(buffer[98]), .B(n419), .C(buffer[97]), .D(n443), .Y(n675)
         );
  INVX1 U773 ( .A(parallel_in[98]), .Y(n674) );
  OAI21X1 U774 ( .A(n368), .B(n676), .C(n677), .Y(n1345) );
  AOI22X1 U775 ( .A(buffer[99]), .B(n419), .C(buffer[98]), .D(n443), .Y(n677)
         );
  INVX1 U776 ( .A(parallel_in[99]), .Y(n676) );
  OAI21X1 U777 ( .A(n368), .B(n678), .C(n679), .Y(n1344) );
  AOI22X1 U778 ( .A(buffer[100]), .B(n418), .C(buffer[99]), .D(n443), .Y(n679)
         );
  INVX1 U779 ( .A(parallel_in[100]), .Y(n678) );
  OAI21X1 U780 ( .A(n368), .B(n680), .C(n681), .Y(n1343) );
  AOI22X1 U781 ( .A(buffer[101]), .B(n418), .C(buffer[100]), .D(n443), .Y(n681) );
  INVX1 U782 ( .A(parallel_in[101]), .Y(n680) );
  OAI21X1 U783 ( .A(n368), .B(n682), .C(n683), .Y(n1342) );
  AOI22X1 U784 ( .A(buffer[102]), .B(n418), .C(buffer[101]), .D(n443), .Y(n683) );
  INVX1 U785 ( .A(parallel_in[102]), .Y(n682) );
  OAI21X1 U786 ( .A(n368), .B(n684), .C(n685), .Y(n1341) );
  AOI22X1 U787 ( .A(buffer[103]), .B(n418), .C(buffer[102]), .D(n443), .Y(n685) );
  INVX1 U788 ( .A(parallel_in[103]), .Y(n684) );
  OAI21X1 U789 ( .A(n369), .B(n686), .C(n687), .Y(n1340) );
  AOI22X1 U790 ( .A(buffer[104]), .B(n418), .C(buffer[103]), .D(n442), .Y(n687) );
  INVX1 U791 ( .A(parallel_in[104]), .Y(n686) );
  OAI21X1 U792 ( .A(n369), .B(n688), .C(n689), .Y(n1339) );
  AOI22X1 U793 ( .A(buffer[105]), .B(n418), .C(buffer[104]), .D(n442), .Y(n689) );
  INVX1 U794 ( .A(parallel_in[105]), .Y(n688) );
  OAI21X1 U795 ( .A(n369), .B(n690), .C(n691), .Y(n1338) );
  AOI22X1 U796 ( .A(buffer[106]), .B(n418), .C(buffer[105]), .D(n442), .Y(n691) );
  INVX1 U797 ( .A(parallel_in[106]), .Y(n690) );
  OAI21X1 U798 ( .A(n369), .B(n692), .C(n693), .Y(n1337) );
  AOI22X1 U799 ( .A(buffer[107]), .B(n418), .C(buffer[106]), .D(n442), .Y(n693) );
  INVX1 U800 ( .A(parallel_in[107]), .Y(n692) );
  OAI21X1 U801 ( .A(n369), .B(n694), .C(n695), .Y(n1336) );
  AOI22X1 U802 ( .A(buffer[108]), .B(n418), .C(buffer[107]), .D(n442), .Y(n695) );
  INVX1 U803 ( .A(parallel_in[108]), .Y(n694) );
  OAI21X1 U804 ( .A(n369), .B(n696), .C(n697), .Y(n1335) );
  AOI22X1 U805 ( .A(buffer[109]), .B(n418), .C(buffer[108]), .D(n442), .Y(n697) );
  INVX1 U806 ( .A(parallel_in[109]), .Y(n696) );
  OAI21X1 U807 ( .A(n369), .B(n698), .C(n699), .Y(n1334) );
  AOI22X1 U808 ( .A(buffer[110]), .B(n418), .C(buffer[109]), .D(n442), .Y(n699) );
  INVX1 U809 ( .A(parallel_in[110]), .Y(n698) );
  OAI21X1 U810 ( .A(n369), .B(n700), .C(n701), .Y(n1333) );
  AOI22X1 U811 ( .A(buffer[111]), .B(n418), .C(buffer[110]), .D(n442), .Y(n701) );
  INVX1 U812 ( .A(parallel_in[111]), .Y(n700) );
  OAI21X1 U813 ( .A(n369), .B(n702), .C(n703), .Y(n1332) );
  AOI22X1 U814 ( .A(buffer[112]), .B(n418), .C(buffer[111]), .D(n442), .Y(n703) );
  INVX1 U815 ( .A(parallel_in[112]), .Y(n702) );
  OAI21X1 U816 ( .A(n369), .B(n704), .C(n705), .Y(n1331) );
  AOI22X1 U817 ( .A(buffer[113]), .B(n417), .C(buffer[112]), .D(n442), .Y(n705) );
  INVX1 U818 ( .A(parallel_in[113]), .Y(n704) );
  OAI21X1 U819 ( .A(n369), .B(n706), .C(n707), .Y(n1330) );
  AOI22X1 U820 ( .A(buffer[114]), .B(n417), .C(buffer[113]), .D(n442), .Y(n707) );
  INVX1 U821 ( .A(parallel_in[114]), .Y(n706) );
  OAI21X1 U822 ( .A(n369), .B(n708), .C(n709), .Y(n1329) );
  AOI22X1 U823 ( .A(buffer[115]), .B(n417), .C(buffer[114]), .D(n442), .Y(n709) );
  INVX1 U824 ( .A(parallel_in[115]), .Y(n708) );
  OAI21X1 U825 ( .A(n369), .B(n710), .C(n711), .Y(n1328) );
  AOI22X1 U826 ( .A(buffer[116]), .B(n417), .C(buffer[115]), .D(n442), .Y(n711) );
  INVX1 U827 ( .A(parallel_in[116]), .Y(n710) );
  OAI21X1 U828 ( .A(n370), .B(n712), .C(n713), .Y(n1327) );
  AOI22X1 U829 ( .A(buffer[117]), .B(n417), .C(buffer[116]), .D(n441), .Y(n713) );
  INVX1 U830 ( .A(parallel_in[117]), .Y(n712) );
  OAI21X1 U831 ( .A(n370), .B(n714), .C(n715), .Y(n1326) );
  AOI22X1 U832 ( .A(buffer[118]), .B(n417), .C(buffer[117]), .D(n441), .Y(n715) );
  INVX1 U833 ( .A(parallel_in[118]), .Y(n714) );
  OAI21X1 U834 ( .A(n370), .B(n716), .C(n717), .Y(n1325) );
  AOI22X1 U835 ( .A(buffer[119]), .B(n417), .C(buffer[118]), .D(n441), .Y(n717) );
  INVX1 U836 ( .A(parallel_in[119]), .Y(n716) );
  OAI21X1 U837 ( .A(n370), .B(n718), .C(n719), .Y(n1324) );
  AOI22X1 U838 ( .A(buffer[120]), .B(n417), .C(buffer[119]), .D(n441), .Y(n719) );
  INVX1 U839 ( .A(parallel_in[120]), .Y(n718) );
  OAI21X1 U840 ( .A(n370), .B(n720), .C(n721), .Y(n1323) );
  AOI22X1 U841 ( .A(buffer[121]), .B(n417), .C(buffer[120]), .D(n441), .Y(n721) );
  INVX1 U842 ( .A(parallel_in[121]), .Y(n720) );
  OAI21X1 U843 ( .A(n370), .B(n722), .C(n723), .Y(n1322) );
  AOI22X1 U844 ( .A(buffer[122]), .B(n417), .C(buffer[121]), .D(n441), .Y(n723) );
  INVX1 U845 ( .A(parallel_in[122]), .Y(n722) );
  OAI21X1 U846 ( .A(n370), .B(n724), .C(n725), .Y(n1321) );
  AOI22X1 U847 ( .A(buffer[123]), .B(n417), .C(buffer[122]), .D(n441), .Y(n725) );
  INVX1 U848 ( .A(parallel_in[123]), .Y(n724) );
  OAI21X1 U849 ( .A(n370), .B(n726), .C(n727), .Y(n1320) );
  AOI22X1 U850 ( .A(buffer[124]), .B(n417), .C(buffer[123]), .D(n441), .Y(n727) );
  INVX1 U851 ( .A(parallel_in[124]), .Y(n726) );
  OAI21X1 U852 ( .A(n370), .B(n728), .C(n729), .Y(n1319) );
  AOI22X1 U853 ( .A(buffer[125]), .B(n417), .C(buffer[124]), .D(n441), .Y(n729) );
  INVX1 U854 ( .A(parallel_in[125]), .Y(n728) );
  OAI21X1 U855 ( .A(n370), .B(n730), .C(n731), .Y(n1318) );
  AOI22X1 U856 ( .A(buffer[126]), .B(n416), .C(buffer[125]), .D(n441), .Y(n731) );
  INVX1 U857 ( .A(parallel_in[126]), .Y(n730) );
  OAI21X1 U858 ( .A(n370), .B(n732), .C(n733), .Y(n1317) );
  AOI22X1 U859 ( .A(buffer[127]), .B(n416), .C(buffer[126]), .D(n441), .Y(n733) );
  INVX1 U860 ( .A(parallel_in[127]), .Y(n732) );
  OAI21X1 U861 ( .A(n370), .B(n734), .C(n735), .Y(n1316) );
  AOI22X1 U862 ( .A(buffer[128]), .B(n416), .C(buffer[127]), .D(n441), .Y(n735) );
  INVX1 U863 ( .A(parallel_in[128]), .Y(n734) );
  OAI21X1 U864 ( .A(n370), .B(n736), .C(n737), .Y(n1315) );
  AOI22X1 U865 ( .A(buffer[129]), .B(n416), .C(buffer[128]), .D(n441), .Y(n737) );
  INVX1 U866 ( .A(parallel_in[129]), .Y(n736) );
  OAI21X1 U867 ( .A(n371), .B(n738), .C(n739), .Y(n1314) );
  AOI22X1 U868 ( .A(buffer[130]), .B(n416), .C(buffer[129]), .D(n440), .Y(n739) );
  INVX1 U869 ( .A(parallel_in[130]), .Y(n738) );
  OAI21X1 U870 ( .A(n371), .B(n740), .C(n741), .Y(n1313) );
  AOI22X1 U871 ( .A(buffer[131]), .B(n416), .C(buffer[130]), .D(n440), .Y(n741) );
  INVX1 U872 ( .A(parallel_in[131]), .Y(n740) );
  OAI21X1 U873 ( .A(n371), .B(n742), .C(n743), .Y(n1312) );
  AOI22X1 U874 ( .A(buffer[132]), .B(n416), .C(buffer[131]), .D(n440), .Y(n743) );
  INVX1 U875 ( .A(parallel_in[132]), .Y(n742) );
  OAI21X1 U876 ( .A(n371), .B(n744), .C(n745), .Y(n1311) );
  AOI22X1 U877 ( .A(buffer[133]), .B(n416), .C(buffer[132]), .D(n440), .Y(n745) );
  INVX1 U878 ( .A(parallel_in[133]), .Y(n744) );
  OAI21X1 U879 ( .A(n371), .B(n746), .C(n747), .Y(n1310) );
  AOI22X1 U880 ( .A(buffer[134]), .B(n416), .C(buffer[133]), .D(n440), .Y(n747) );
  INVX1 U881 ( .A(parallel_in[134]), .Y(n746) );
  OAI21X1 U882 ( .A(n371), .B(n748), .C(n749), .Y(n1309) );
  AOI22X1 U883 ( .A(buffer[135]), .B(n416), .C(buffer[134]), .D(n440), .Y(n749) );
  INVX1 U884 ( .A(parallel_in[135]), .Y(n748) );
  OAI21X1 U885 ( .A(n371), .B(n750), .C(n751), .Y(n1308) );
  AOI22X1 U886 ( .A(buffer[136]), .B(n416), .C(buffer[135]), .D(n440), .Y(n751) );
  INVX1 U887 ( .A(parallel_in[136]), .Y(n750) );
  OAI21X1 U888 ( .A(n371), .B(n752), .C(n753), .Y(n1307) );
  AOI22X1 U889 ( .A(buffer[137]), .B(n416), .C(buffer[136]), .D(n440), .Y(n753) );
  INVX1 U890 ( .A(parallel_in[137]), .Y(n752) );
  OAI21X1 U891 ( .A(n371), .B(n754), .C(n755), .Y(n1306) );
  AOI22X1 U892 ( .A(buffer[138]), .B(n416), .C(buffer[137]), .D(n440), .Y(n755) );
  INVX1 U893 ( .A(parallel_in[138]), .Y(n754) );
  OAI21X1 U894 ( .A(n371), .B(n756), .C(n757), .Y(n1305) );
  AOI22X1 U895 ( .A(buffer[139]), .B(n415), .C(buffer[138]), .D(n440), .Y(n757) );
  INVX1 U896 ( .A(parallel_in[139]), .Y(n756) );
  OAI21X1 U897 ( .A(n371), .B(n758), .C(n759), .Y(n1304) );
  AOI22X1 U898 ( .A(buffer[140]), .B(n415), .C(buffer[139]), .D(n440), .Y(n759) );
  INVX1 U899 ( .A(parallel_in[140]), .Y(n758) );
  OAI21X1 U900 ( .A(n371), .B(n760), .C(n761), .Y(n1303) );
  AOI22X1 U901 ( .A(buffer[141]), .B(n415), .C(buffer[140]), .D(n440), .Y(n761) );
  INVX1 U902 ( .A(parallel_in[141]), .Y(n760) );
  OAI21X1 U903 ( .A(n371), .B(n762), .C(n763), .Y(n1302) );
  AOI22X1 U904 ( .A(buffer[142]), .B(n415), .C(buffer[141]), .D(n440), .Y(n763) );
  INVX1 U905 ( .A(parallel_in[142]), .Y(n762) );
  OAI21X1 U906 ( .A(n372), .B(n764), .C(n765), .Y(n1301) );
  AOI22X1 U907 ( .A(buffer[143]), .B(n415), .C(buffer[142]), .D(n439), .Y(n765) );
  INVX1 U908 ( .A(parallel_in[143]), .Y(n764) );
  OAI21X1 U909 ( .A(n372), .B(n766), .C(n767), .Y(n1300) );
  AOI22X1 U910 ( .A(buffer[144]), .B(n415), .C(buffer[143]), .D(n439), .Y(n767) );
  INVX1 U911 ( .A(parallel_in[144]), .Y(n766) );
  OAI21X1 U912 ( .A(n372), .B(n768), .C(n769), .Y(n1299) );
  AOI22X1 U913 ( .A(buffer[145]), .B(n415), .C(buffer[144]), .D(n439), .Y(n769) );
  INVX1 U914 ( .A(parallel_in[145]), .Y(n768) );
  OAI21X1 U915 ( .A(n372), .B(n770), .C(n771), .Y(n1298) );
  AOI22X1 U916 ( .A(buffer[146]), .B(n415), .C(buffer[145]), .D(n439), .Y(n771) );
  INVX1 U917 ( .A(parallel_in[146]), .Y(n770) );
  OAI21X1 U918 ( .A(n372), .B(n772), .C(n773), .Y(n1297) );
  AOI22X1 U919 ( .A(buffer[147]), .B(n415), .C(buffer[146]), .D(n439), .Y(n773) );
  INVX1 U920 ( .A(parallel_in[147]), .Y(n772) );
  OAI21X1 U921 ( .A(n372), .B(n774), .C(n775), .Y(n1296) );
  AOI22X1 U922 ( .A(buffer[148]), .B(n415), .C(buffer[147]), .D(n439), .Y(n775) );
  INVX1 U923 ( .A(parallel_in[148]), .Y(n774) );
  OAI21X1 U924 ( .A(n372), .B(n776), .C(n777), .Y(n1295) );
  AOI22X1 U925 ( .A(buffer[149]), .B(n415), .C(buffer[148]), .D(n439), .Y(n777) );
  INVX1 U926 ( .A(parallel_in[149]), .Y(n776) );
  OAI21X1 U927 ( .A(n372), .B(n778), .C(n779), .Y(n1294) );
  AOI22X1 U928 ( .A(buffer[150]), .B(n415), .C(buffer[149]), .D(n439), .Y(n779) );
  INVX1 U929 ( .A(parallel_in[150]), .Y(n778) );
  OAI21X1 U930 ( .A(n372), .B(n780), .C(n781), .Y(n1293) );
  AOI22X1 U931 ( .A(buffer[151]), .B(n415), .C(buffer[150]), .D(n439), .Y(n781) );
  INVX1 U932 ( .A(parallel_in[151]), .Y(n780) );
  OAI21X1 U933 ( .A(n372), .B(n782), .C(n783), .Y(n1292) );
  AOI22X1 U934 ( .A(buffer[152]), .B(n414), .C(buffer[151]), .D(n439), .Y(n783) );
  INVX1 U935 ( .A(parallel_in[152]), .Y(n782) );
  OAI21X1 U936 ( .A(n372), .B(n784), .C(n785), .Y(n1291) );
  AOI22X1 U937 ( .A(buffer[153]), .B(n414), .C(buffer[152]), .D(n439), .Y(n785) );
  INVX1 U938 ( .A(parallel_in[153]), .Y(n784) );
  OAI21X1 U939 ( .A(n372), .B(n786), .C(n787), .Y(n1290) );
  AOI22X1 U940 ( .A(buffer[154]), .B(n414), .C(buffer[153]), .D(n439), .Y(n787) );
  INVX1 U941 ( .A(parallel_in[154]), .Y(n786) );
  OAI21X1 U942 ( .A(n372), .B(n788), .C(n789), .Y(n1289) );
  AOI22X1 U943 ( .A(buffer[155]), .B(n414), .C(buffer[154]), .D(n439), .Y(n789) );
  INVX1 U944 ( .A(parallel_in[155]), .Y(n788) );
  OAI21X1 U945 ( .A(n373), .B(n790), .C(n791), .Y(n1288) );
  AOI22X1 U946 ( .A(buffer[156]), .B(n414), .C(buffer[155]), .D(n438), .Y(n791) );
  INVX1 U947 ( .A(parallel_in[156]), .Y(n790) );
  OAI21X1 U948 ( .A(n373), .B(n792), .C(n793), .Y(n1287) );
  AOI22X1 U949 ( .A(buffer[157]), .B(n414), .C(buffer[156]), .D(n438), .Y(n793) );
  INVX1 U950 ( .A(parallel_in[157]), .Y(n792) );
  OAI21X1 U951 ( .A(n373), .B(n794), .C(n795), .Y(n1286) );
  AOI22X1 U952 ( .A(buffer[158]), .B(n414), .C(buffer[157]), .D(n438), .Y(n795) );
  INVX1 U953 ( .A(parallel_in[158]), .Y(n794) );
  OAI21X1 U954 ( .A(n373), .B(n796), .C(n797), .Y(n1285) );
  AOI22X1 U955 ( .A(buffer[159]), .B(n414), .C(buffer[158]), .D(n438), .Y(n797) );
  INVX1 U956 ( .A(parallel_in[159]), .Y(n796) );
  OAI21X1 U957 ( .A(n373), .B(n798), .C(n799), .Y(n1284) );
  AOI22X1 U958 ( .A(buffer[160]), .B(n414), .C(buffer[159]), .D(n438), .Y(n799) );
  INVX1 U959 ( .A(parallel_in[160]), .Y(n798) );
  OAI21X1 U960 ( .A(n373), .B(n800), .C(n801), .Y(n1283) );
  AOI22X1 U961 ( .A(buffer[161]), .B(n414), .C(buffer[160]), .D(n438), .Y(n801) );
  INVX1 U962 ( .A(parallel_in[161]), .Y(n800) );
  OAI21X1 U963 ( .A(n373), .B(n802), .C(n803), .Y(n1282) );
  AOI22X1 U964 ( .A(buffer[162]), .B(n414), .C(buffer[161]), .D(n438), .Y(n803) );
  INVX1 U965 ( .A(parallel_in[162]), .Y(n802) );
  OAI21X1 U966 ( .A(n373), .B(n804), .C(n805), .Y(n1281) );
  AOI22X1 U967 ( .A(buffer[163]), .B(n414), .C(buffer[162]), .D(n438), .Y(n805) );
  INVX1 U968 ( .A(parallel_in[163]), .Y(n804) );
  OAI21X1 U969 ( .A(n373), .B(n806), .C(n807), .Y(n1280) );
  AOI22X1 U970 ( .A(buffer[164]), .B(n414), .C(buffer[163]), .D(n438), .Y(n807) );
  INVX1 U971 ( .A(parallel_in[164]), .Y(n806) );
  OAI21X1 U972 ( .A(n373), .B(n808), .C(n809), .Y(n1279) );
  AOI22X1 U973 ( .A(buffer[165]), .B(n413), .C(buffer[164]), .D(n438), .Y(n809) );
  INVX1 U974 ( .A(parallel_in[165]), .Y(n808) );
  OAI21X1 U975 ( .A(n373), .B(n810), .C(n811), .Y(n1278) );
  AOI22X1 U976 ( .A(buffer[166]), .B(n413), .C(buffer[165]), .D(n438), .Y(n811) );
  INVX1 U977 ( .A(parallel_in[166]), .Y(n810) );
  OAI21X1 U978 ( .A(n373), .B(n812), .C(n813), .Y(n1277) );
  AOI22X1 U979 ( .A(buffer[167]), .B(n413), .C(buffer[166]), .D(n438), .Y(n813) );
  INVX1 U980 ( .A(parallel_in[167]), .Y(n812) );
  OAI21X1 U981 ( .A(n373), .B(n814), .C(n815), .Y(n1276) );
  AOI22X1 U982 ( .A(buffer[168]), .B(n413), .C(buffer[167]), .D(n438), .Y(n815) );
  INVX1 U983 ( .A(parallel_in[168]), .Y(n814) );
  OAI21X1 U984 ( .A(n374), .B(n816), .C(n817), .Y(n1275) );
  AOI22X1 U985 ( .A(buffer[169]), .B(n413), .C(buffer[168]), .D(n437), .Y(n817) );
  INVX1 U986 ( .A(parallel_in[169]), .Y(n816) );
  OAI21X1 U987 ( .A(n374), .B(n818), .C(n819), .Y(n1274) );
  AOI22X1 U988 ( .A(buffer[170]), .B(n413), .C(buffer[169]), .D(n437), .Y(n819) );
  INVX1 U989 ( .A(parallel_in[170]), .Y(n818) );
  OAI21X1 U990 ( .A(n374), .B(n820), .C(n821), .Y(n1273) );
  AOI22X1 U991 ( .A(buffer[171]), .B(n413), .C(buffer[170]), .D(n437), .Y(n821) );
  INVX1 U992 ( .A(parallel_in[171]), .Y(n820) );
  OAI21X1 U993 ( .A(n374), .B(n822), .C(n823), .Y(n1272) );
  AOI22X1 U994 ( .A(buffer[172]), .B(n413), .C(buffer[171]), .D(n437), .Y(n823) );
  INVX1 U995 ( .A(parallel_in[172]), .Y(n822) );
  OAI21X1 U996 ( .A(n374), .B(n824), .C(n825), .Y(n1271) );
  AOI22X1 U997 ( .A(buffer[173]), .B(n413), .C(buffer[172]), .D(n437), .Y(n825) );
  INVX1 U998 ( .A(parallel_in[173]), .Y(n824) );
  OAI21X1 U999 ( .A(n374), .B(n826), .C(n827), .Y(n1270) );
  AOI22X1 U1000 ( .A(buffer[174]), .B(n413), .C(buffer[173]), .D(n437), .Y(
        n827) );
  INVX1 U1001 ( .A(parallel_in[174]), .Y(n826) );
  OAI21X1 U1002 ( .A(n374), .B(n828), .C(n829), .Y(n1269) );
  AOI22X1 U1003 ( .A(buffer[175]), .B(n413), .C(buffer[174]), .D(n437), .Y(
        n829) );
  INVX1 U1004 ( .A(parallel_in[175]), .Y(n828) );
  OAI21X1 U1005 ( .A(n374), .B(n830), .C(n831), .Y(n1268) );
  AOI22X1 U1006 ( .A(buffer[176]), .B(n413), .C(buffer[175]), .D(n437), .Y(
        n831) );
  INVX1 U1007 ( .A(parallel_in[176]), .Y(n830) );
  OAI21X1 U1008 ( .A(n374), .B(n832), .C(n833), .Y(n1267) );
  AOI22X1 U1009 ( .A(buffer[177]), .B(n413), .C(buffer[176]), .D(n437), .Y(
        n833) );
  INVX1 U1010 ( .A(parallel_in[177]), .Y(n832) );
  OAI21X1 U1011 ( .A(n374), .B(n834), .C(n835), .Y(n1266) );
  AOI22X1 U1012 ( .A(buffer[178]), .B(n412), .C(buffer[177]), .D(n437), .Y(
        n835) );
  INVX1 U1013 ( .A(parallel_in[178]), .Y(n834) );
  OAI21X1 U1014 ( .A(n374), .B(n836), .C(n837), .Y(n1265) );
  AOI22X1 U1015 ( .A(buffer[179]), .B(n412), .C(buffer[178]), .D(n437), .Y(
        n837) );
  INVX1 U1016 ( .A(parallel_in[179]), .Y(n836) );
  OAI21X1 U1017 ( .A(n374), .B(n838), .C(n839), .Y(n1264) );
  AOI22X1 U1018 ( .A(buffer[180]), .B(n412), .C(buffer[179]), .D(n437), .Y(
        n839) );
  INVX1 U1019 ( .A(parallel_in[180]), .Y(n838) );
  OAI21X1 U1020 ( .A(n374), .B(n840), .C(n841), .Y(n1263) );
  AOI22X1 U1021 ( .A(buffer[181]), .B(n412), .C(buffer[180]), .D(n443), .Y(
        n841) );
  INVX1 U1022 ( .A(parallel_in[181]), .Y(n840) );
  OAI21X1 U1023 ( .A(n375), .B(n842), .C(n843), .Y(n1262) );
  AOI22X1 U1024 ( .A(buffer[182]), .B(n412), .C(buffer[181]), .D(n464), .Y(
        n843) );
  INVX1 U1025 ( .A(parallel_in[182]), .Y(n842) );
  OAI21X1 U1026 ( .A(n375), .B(n844), .C(n845), .Y(n1261) );
  AOI22X1 U1027 ( .A(buffer[183]), .B(n412), .C(buffer[182]), .D(n464), .Y(
        n845) );
  INVX1 U1028 ( .A(parallel_in[183]), .Y(n844) );
  OAI21X1 U1029 ( .A(n375), .B(n846), .C(n847), .Y(n1260) );
  AOI22X1 U1030 ( .A(buffer[184]), .B(n412), .C(buffer[183]), .D(n464), .Y(
        n847) );
  INVX1 U1031 ( .A(parallel_in[184]), .Y(n846) );
  OAI21X1 U1032 ( .A(n375), .B(n848), .C(n849), .Y(n1259) );
  AOI22X1 U1033 ( .A(buffer[185]), .B(n412), .C(buffer[184]), .D(n464), .Y(
        n849) );
  INVX1 U1034 ( .A(parallel_in[185]), .Y(n848) );
  OAI21X1 U1035 ( .A(n375), .B(n850), .C(n851), .Y(n1258) );
  AOI22X1 U1036 ( .A(buffer[186]), .B(n412), .C(buffer[185]), .D(n463), .Y(
        n851) );
  INVX1 U1037 ( .A(parallel_in[186]), .Y(n850) );
  OAI21X1 U1038 ( .A(n375), .B(n852), .C(n853), .Y(n1257) );
  AOI22X1 U1039 ( .A(buffer[187]), .B(n412), .C(buffer[186]), .D(n464), .Y(
        n853) );
  INVX1 U1040 ( .A(parallel_in[187]), .Y(n852) );
  OAI21X1 U1041 ( .A(n375), .B(n854), .C(n855), .Y(n1256) );
  AOI22X1 U1042 ( .A(buffer[188]), .B(n412), .C(buffer[187]), .D(n464), .Y(
        n855) );
  INVX1 U1043 ( .A(parallel_in[188]), .Y(n854) );
  OAI21X1 U1044 ( .A(n375), .B(n856), .C(n857), .Y(n1255) );
  AOI22X1 U1045 ( .A(buffer[189]), .B(n412), .C(buffer[188]), .D(n463), .Y(
        n857) );
  INVX1 U1046 ( .A(parallel_in[189]), .Y(n856) );
  OAI21X1 U1047 ( .A(n375), .B(n858), .C(n859), .Y(n1254) );
  AOI22X1 U1048 ( .A(buffer[190]), .B(n412), .C(buffer[189]), .D(n463), .Y(
        n859) );
  INVX1 U1049 ( .A(parallel_in[190]), .Y(n858) );
  OAI21X1 U1050 ( .A(n375), .B(n860), .C(n861), .Y(n1253) );
  AOI22X1 U1051 ( .A(buffer[191]), .B(n411), .C(buffer[190]), .D(n463), .Y(
        n861) );
  INVX1 U1052 ( .A(parallel_in[191]), .Y(n860) );
  OAI21X1 U1053 ( .A(n375), .B(n862), .C(n863), .Y(n1252) );
  AOI22X1 U1054 ( .A(buffer[192]), .B(n411), .C(buffer[191]), .D(n463), .Y(
        n863) );
  INVX1 U1055 ( .A(parallel_in[192]), .Y(n862) );
  OAI21X1 U1056 ( .A(n375), .B(n864), .C(n865), .Y(n1251) );
  AOI22X1 U1057 ( .A(buffer[193]), .B(n411), .C(buffer[192]), .D(n463), .Y(
        n865) );
  INVX1 U1058 ( .A(parallel_in[193]), .Y(n864) );
  OAI21X1 U1059 ( .A(n375), .B(n866), .C(n867), .Y(n1250) );
  AOI22X1 U1060 ( .A(buffer[194]), .B(n411), .C(buffer[193]), .D(n463), .Y(
        n867) );
  INVX1 U1061 ( .A(parallel_in[194]), .Y(n866) );
  OAI21X1 U1062 ( .A(n376), .B(n868), .C(n869), .Y(n1249) );
  AOI22X1 U1063 ( .A(buffer[195]), .B(n411), .C(buffer[194]), .D(n463), .Y(
        n869) );
  INVX1 U1064 ( .A(parallel_in[195]), .Y(n868) );
  OAI21X1 U1065 ( .A(n376), .B(n870), .C(n871), .Y(n1248) );
  AOI22X1 U1066 ( .A(buffer[196]), .B(n411), .C(buffer[195]), .D(n463), .Y(
        n871) );
  INVX1 U1067 ( .A(parallel_in[196]), .Y(n870) );
  OAI21X1 U1068 ( .A(n376), .B(n872), .C(n873), .Y(n1247) );
  AOI22X1 U1069 ( .A(buffer[197]), .B(n411), .C(buffer[196]), .D(n463), .Y(
        n873) );
  INVX1 U1070 ( .A(parallel_in[197]), .Y(n872) );
  OAI21X1 U1071 ( .A(n376), .B(n874), .C(n875), .Y(n1246) );
  AOI22X1 U1072 ( .A(buffer[198]), .B(n411), .C(buffer[197]), .D(n463), .Y(
        n875) );
  INVX1 U1073 ( .A(parallel_in[198]), .Y(n874) );
  OAI21X1 U1074 ( .A(n376), .B(n876), .C(n877), .Y(n1245) );
  AOI22X1 U1075 ( .A(buffer[199]), .B(n411), .C(buffer[198]), .D(n463), .Y(
        n877) );
  INVX1 U1076 ( .A(parallel_in[199]), .Y(n876) );
  OAI21X1 U1077 ( .A(n376), .B(n878), .C(n879), .Y(n1244) );
  AOI22X1 U1078 ( .A(buffer[200]), .B(n411), .C(buffer[199]), .D(n463), .Y(
        n879) );
  INVX1 U1079 ( .A(parallel_in[200]), .Y(n878) );
  OAI21X1 U1080 ( .A(n376), .B(n880), .C(n881), .Y(n1243) );
  AOI22X1 U1081 ( .A(buffer[201]), .B(n411), .C(buffer[200]), .D(n462), .Y(
        n881) );
  INVX1 U1082 ( .A(parallel_in[201]), .Y(n880) );
  OAI21X1 U1083 ( .A(n376), .B(n882), .C(n883), .Y(n1242) );
  AOI22X1 U1084 ( .A(buffer[202]), .B(n411), .C(buffer[201]), .D(n462), .Y(
        n883) );
  INVX1 U1085 ( .A(parallel_in[202]), .Y(n882) );
  OAI21X1 U1086 ( .A(n376), .B(n884), .C(n885), .Y(n1241) );
  AOI22X1 U1087 ( .A(buffer[203]), .B(n411), .C(buffer[202]), .D(n462), .Y(
        n885) );
  INVX1 U1088 ( .A(parallel_in[203]), .Y(n884) );
  OAI21X1 U1089 ( .A(n376), .B(n886), .C(n887), .Y(n1240) );
  AOI22X1 U1090 ( .A(buffer[204]), .B(n410), .C(buffer[203]), .D(n462), .Y(
        n887) );
  INVX1 U1091 ( .A(parallel_in[204]), .Y(n886) );
  OAI21X1 U1092 ( .A(n376), .B(n888), .C(n889), .Y(n1239) );
  AOI22X1 U1093 ( .A(buffer[205]), .B(n410), .C(buffer[204]), .D(n462), .Y(
        n889) );
  INVX1 U1094 ( .A(parallel_in[205]), .Y(n888) );
  OAI21X1 U1095 ( .A(n376), .B(n890), .C(n891), .Y(n1238) );
  AOI22X1 U1096 ( .A(buffer[206]), .B(n410), .C(buffer[205]), .D(n462), .Y(
        n891) );
  INVX1 U1097 ( .A(parallel_in[206]), .Y(n890) );
  OAI21X1 U1098 ( .A(n376), .B(n892), .C(n893), .Y(n1237) );
  AOI22X1 U1099 ( .A(buffer[207]), .B(n410), .C(buffer[206]), .D(n462), .Y(
        n893) );
  INVX1 U1100 ( .A(parallel_in[207]), .Y(n892) );
  OAI21X1 U1101 ( .A(n377), .B(n894), .C(n895), .Y(n1236) );
  AOI22X1 U1102 ( .A(buffer[208]), .B(n410), .C(buffer[207]), .D(n462), .Y(
        n895) );
  INVX1 U1103 ( .A(parallel_in[208]), .Y(n894) );
  OAI21X1 U1104 ( .A(n377), .B(n896), .C(n897), .Y(n1235) );
  AOI22X1 U1105 ( .A(buffer[209]), .B(n410), .C(buffer[208]), .D(n462), .Y(
        n897) );
  INVX1 U1106 ( .A(parallel_in[209]), .Y(n896) );
  OAI21X1 U1107 ( .A(n377), .B(n898), .C(n899), .Y(n1234) );
  AOI22X1 U1108 ( .A(buffer[210]), .B(n410), .C(buffer[209]), .D(n462), .Y(
        n899) );
  INVX1 U1109 ( .A(parallel_in[210]), .Y(n898) );
  OAI21X1 U1110 ( .A(n377), .B(n900), .C(n901), .Y(n1233) );
  AOI22X1 U1111 ( .A(buffer[211]), .B(n410), .C(buffer[210]), .D(n462), .Y(
        n901) );
  INVX1 U1112 ( .A(parallel_in[211]), .Y(n900) );
  OAI21X1 U1113 ( .A(n377), .B(n902), .C(n903), .Y(n1232) );
  AOI22X1 U1114 ( .A(buffer[212]), .B(n410), .C(buffer[211]), .D(n462), .Y(
        n903) );
  INVX1 U1115 ( .A(parallel_in[212]), .Y(n902) );
  OAI21X1 U1116 ( .A(n377), .B(n904), .C(n905), .Y(n1231) );
  AOI22X1 U1117 ( .A(buffer[213]), .B(n410), .C(buffer[212]), .D(n461), .Y(
        n905) );
  INVX1 U1118 ( .A(parallel_in[213]), .Y(n904) );
  OAI21X1 U1119 ( .A(n377), .B(n906), .C(n907), .Y(n1230) );
  AOI22X1 U1120 ( .A(buffer[214]), .B(n410), .C(buffer[213]), .D(n462), .Y(
        n907) );
  INVX1 U1121 ( .A(parallel_in[214]), .Y(n906) );
  OAI21X1 U1122 ( .A(n377), .B(n908), .C(n909), .Y(n1229) );
  AOI22X1 U1123 ( .A(buffer[215]), .B(n410), .C(buffer[214]), .D(n461), .Y(
        n909) );
  INVX1 U1124 ( .A(parallel_in[215]), .Y(n908) );
  OAI21X1 U1125 ( .A(n377), .B(n910), .C(n911), .Y(n1228) );
  AOI22X1 U1126 ( .A(buffer[216]), .B(n410), .C(buffer[215]), .D(n461), .Y(
        n911) );
  INVX1 U1127 ( .A(parallel_in[216]), .Y(n910) );
  OAI21X1 U1128 ( .A(n377), .B(n912), .C(n913), .Y(n1227) );
  AOI22X1 U1129 ( .A(buffer[217]), .B(n409), .C(buffer[216]), .D(n461), .Y(
        n913) );
  INVX1 U1130 ( .A(parallel_in[217]), .Y(n912) );
  OAI21X1 U1131 ( .A(n377), .B(n914), .C(n915), .Y(n1226) );
  AOI22X1 U1132 ( .A(buffer[218]), .B(n409), .C(buffer[217]), .D(n461), .Y(
        n915) );
  INVX1 U1133 ( .A(parallel_in[218]), .Y(n914) );
  OAI21X1 U1134 ( .A(n377), .B(n916), .C(n917), .Y(n1225) );
  AOI22X1 U1135 ( .A(buffer[219]), .B(n409), .C(buffer[218]), .D(n461), .Y(
        n917) );
  INVX1 U1136 ( .A(parallel_in[219]), .Y(n916) );
  OAI21X1 U1137 ( .A(n377), .B(n918), .C(n919), .Y(n1224) );
  AOI22X1 U1138 ( .A(buffer[220]), .B(n409), .C(buffer[219]), .D(n461), .Y(
        n919) );
  INVX1 U1139 ( .A(parallel_in[220]), .Y(n918) );
  OAI21X1 U1140 ( .A(n378), .B(n920), .C(n921), .Y(n1223) );
  AOI22X1 U1141 ( .A(buffer[221]), .B(n409), .C(buffer[220]), .D(n461), .Y(
        n921) );
  INVX1 U1142 ( .A(parallel_in[221]), .Y(n920) );
  OAI21X1 U1143 ( .A(n378), .B(n922), .C(n923), .Y(n1222) );
  AOI22X1 U1144 ( .A(buffer[222]), .B(n409), .C(buffer[221]), .D(n461), .Y(
        n923) );
  INVX1 U1145 ( .A(parallel_in[222]), .Y(n922) );
  OAI21X1 U1146 ( .A(n378), .B(n924), .C(n925), .Y(n1221) );
  AOI22X1 U1147 ( .A(buffer[223]), .B(n409), .C(buffer[222]), .D(n461), .Y(
        n925) );
  INVX1 U1148 ( .A(parallel_in[223]), .Y(n924) );
  OAI21X1 U1149 ( .A(n378), .B(n926), .C(n927), .Y(n1220) );
  AOI22X1 U1150 ( .A(buffer[224]), .B(n409), .C(buffer[223]), .D(n461), .Y(
        n927) );
  INVX1 U1151 ( .A(parallel_in[224]), .Y(n926) );
  OAI21X1 U1152 ( .A(n378), .B(n928), .C(n929), .Y(n1219) );
  AOI22X1 U1153 ( .A(buffer[225]), .B(n409), .C(buffer[224]), .D(n461), .Y(
        n929) );
  INVX1 U1154 ( .A(parallel_in[225]), .Y(n928) );
  OAI21X1 U1155 ( .A(n378), .B(n930), .C(n931), .Y(n1218) );
  AOI22X1 U1156 ( .A(buffer[226]), .B(n409), .C(buffer[225]), .D(n461), .Y(
        n931) );
  INVX1 U1157 ( .A(parallel_in[226]), .Y(n930) );
  OAI21X1 U1158 ( .A(n378), .B(n932), .C(n933), .Y(n1217) );
  AOI22X1 U1159 ( .A(buffer[227]), .B(n409), .C(buffer[226]), .D(n460), .Y(
        n933) );
  INVX1 U1160 ( .A(parallel_in[227]), .Y(n932) );
  OAI21X1 U1161 ( .A(n378), .B(n934), .C(n935), .Y(n1216) );
  AOI22X1 U1162 ( .A(buffer[228]), .B(n409), .C(buffer[227]), .D(n460), .Y(
        n935) );
  INVX1 U1163 ( .A(parallel_in[228]), .Y(n934) );
  OAI21X1 U1164 ( .A(n378), .B(n936), .C(n937), .Y(n1215) );
  AOI22X1 U1165 ( .A(buffer[229]), .B(n409), .C(buffer[228]), .D(n460), .Y(
        n937) );
  INVX1 U1166 ( .A(parallel_in[229]), .Y(n936) );
  OAI21X1 U1167 ( .A(n378), .B(n938), .C(n939), .Y(n1214) );
  AOI22X1 U1168 ( .A(buffer[230]), .B(n408), .C(buffer[229]), .D(n460), .Y(
        n939) );
  INVX1 U1169 ( .A(parallel_in[230]), .Y(n938) );
  OAI21X1 U1170 ( .A(n378), .B(n940), .C(n941), .Y(n1213) );
  AOI22X1 U1171 ( .A(buffer[231]), .B(n408), .C(buffer[230]), .D(n460), .Y(
        n941) );
  INVX1 U1172 ( .A(parallel_in[231]), .Y(n940) );
  OAI21X1 U1173 ( .A(n378), .B(n942), .C(n943), .Y(n1212) );
  AOI22X1 U1174 ( .A(buffer[232]), .B(n408), .C(buffer[231]), .D(n460), .Y(
        n943) );
  INVX1 U1175 ( .A(parallel_in[232]), .Y(n942) );
  OAI21X1 U1176 ( .A(n378), .B(n944), .C(n945), .Y(n1211) );
  AOI22X1 U1177 ( .A(buffer[233]), .B(n408), .C(buffer[232]), .D(n460), .Y(
        n945) );
  INVX1 U1178 ( .A(parallel_in[233]), .Y(n944) );
  OAI21X1 U1179 ( .A(n379), .B(n946), .C(n947), .Y(n1210) );
  AOI22X1 U1180 ( .A(buffer[234]), .B(n408), .C(buffer[233]), .D(n460), .Y(
        n947) );
  INVX1 U1181 ( .A(parallel_in[234]), .Y(n946) );
  OAI21X1 U1182 ( .A(n379), .B(n948), .C(n949), .Y(n1209) );
  AOI22X1 U1183 ( .A(buffer[235]), .B(n408), .C(buffer[234]), .D(n460), .Y(
        n949) );
  INVX1 U1184 ( .A(parallel_in[235]), .Y(n948) );
  OAI21X1 U1185 ( .A(n379), .B(n950), .C(n951), .Y(n1208) );
  AOI22X1 U1186 ( .A(buffer[236]), .B(n408), .C(buffer[235]), .D(n460), .Y(
        n951) );
  INVX1 U1187 ( .A(parallel_in[236]), .Y(n950) );
  OAI21X1 U1188 ( .A(n379), .B(n952), .C(n953), .Y(n1207) );
  AOI22X1 U1189 ( .A(buffer[237]), .B(n408), .C(buffer[236]), .D(n460), .Y(
        n953) );
  INVX1 U1190 ( .A(parallel_in[237]), .Y(n952) );
  OAI21X1 U1191 ( .A(n379), .B(n954), .C(n955), .Y(n1206) );
  AOI22X1 U1192 ( .A(buffer[238]), .B(n408), .C(buffer[237]), .D(n460), .Y(
        n955) );
  INVX1 U1193 ( .A(parallel_in[238]), .Y(n954) );
  OAI21X1 U1194 ( .A(n379), .B(n956), .C(n957), .Y(n1205) );
  AOI22X1 U1195 ( .A(buffer[239]), .B(n408), .C(buffer[238]), .D(n459), .Y(
        n957) );
  INVX1 U1196 ( .A(parallel_in[239]), .Y(n956) );
  OAI21X1 U1197 ( .A(n379), .B(n958), .C(n959), .Y(n1204) );
  AOI22X1 U1198 ( .A(buffer[240]), .B(n408), .C(buffer[239]), .D(n460), .Y(
        n959) );
  INVX1 U1199 ( .A(parallel_in[240]), .Y(n958) );
  OAI21X1 U1200 ( .A(n379), .B(n960), .C(n961), .Y(n1203) );
  AOI22X1 U1201 ( .A(buffer[241]), .B(n408), .C(buffer[240]), .D(n459), .Y(
        n961) );
  INVX1 U1202 ( .A(parallel_in[241]), .Y(n960) );
  OAI21X1 U1203 ( .A(n379), .B(n962), .C(n963), .Y(n1202) );
  AOI22X1 U1204 ( .A(buffer[242]), .B(n408), .C(buffer[241]), .D(n459), .Y(
        n963) );
  INVX1 U1205 ( .A(parallel_in[242]), .Y(n962) );
  OAI21X1 U1206 ( .A(n379), .B(n964), .C(n965), .Y(n1201) );
  AOI22X1 U1207 ( .A(buffer[243]), .B(n407), .C(buffer[242]), .D(n459), .Y(
        n965) );
  INVX1 U1208 ( .A(parallel_in[243]), .Y(n964) );
  OAI21X1 U1209 ( .A(n379), .B(n966), .C(n967), .Y(n1200) );
  AOI22X1 U1210 ( .A(buffer[244]), .B(n407), .C(buffer[243]), .D(n459), .Y(
        n967) );
  INVX1 U1211 ( .A(parallel_in[244]), .Y(n966) );
  OAI21X1 U1212 ( .A(n379), .B(n968), .C(n969), .Y(n1199) );
  AOI22X1 U1213 ( .A(buffer[245]), .B(n407), .C(buffer[244]), .D(n459), .Y(
        n969) );
  INVX1 U1214 ( .A(parallel_in[245]), .Y(n968) );
  OAI21X1 U1215 ( .A(n379), .B(n970), .C(n971), .Y(n1198) );
  AOI22X1 U1216 ( .A(buffer[246]), .B(n407), .C(buffer[245]), .D(n459), .Y(
        n971) );
  INVX1 U1217 ( .A(parallel_in[246]), .Y(n970) );
  OAI21X1 U1218 ( .A(n380), .B(n972), .C(n973), .Y(n1197) );
  AOI22X1 U1219 ( .A(buffer[247]), .B(n407), .C(buffer[246]), .D(n459), .Y(
        n973) );
  INVX1 U1220 ( .A(parallel_in[247]), .Y(n972) );
  OAI21X1 U1221 ( .A(n380), .B(n974), .C(n975), .Y(n1196) );
  AOI22X1 U1222 ( .A(buffer[248]), .B(n407), .C(buffer[247]), .D(n459), .Y(
        n975) );
  INVX1 U1223 ( .A(parallel_in[248]), .Y(n974) );
  OAI21X1 U1224 ( .A(n380), .B(n976), .C(n977), .Y(n1195) );
  AOI22X1 U1225 ( .A(buffer[249]), .B(n407), .C(buffer[248]), .D(n459), .Y(
        n977) );
  INVX1 U1226 ( .A(parallel_in[249]), .Y(n976) );
  OAI21X1 U1227 ( .A(n380), .B(n978), .C(n979), .Y(n1194) );
  AOI22X1 U1228 ( .A(buffer[250]), .B(n407), .C(buffer[249]), .D(n459), .Y(
        n979) );
  INVX1 U1229 ( .A(parallel_in[250]), .Y(n978) );
  OAI21X1 U1230 ( .A(n380), .B(n980), .C(n981), .Y(n1193) );
  AOI22X1 U1231 ( .A(buffer[251]), .B(n407), .C(buffer[250]), .D(n458), .Y(
        n981) );
  INVX1 U1232 ( .A(parallel_in[251]), .Y(n980) );
  OAI21X1 U1233 ( .A(n380), .B(n982), .C(n983), .Y(n1192) );
  AOI22X1 U1234 ( .A(buffer[252]), .B(n407), .C(buffer[251]), .D(n459), .Y(
        n983) );
  INVX1 U1235 ( .A(parallel_in[252]), .Y(n982) );
  OAI21X1 U1236 ( .A(n380), .B(n984), .C(n985), .Y(n1191) );
  AOI22X1 U1237 ( .A(buffer[253]), .B(n407), .C(buffer[252]), .D(n459), .Y(
        n985) );
  INVX1 U1238 ( .A(parallel_in[253]), .Y(n984) );
  OAI21X1 U1239 ( .A(n380), .B(n986), .C(n987), .Y(n1190) );
  AOI22X1 U1240 ( .A(buffer[254]), .B(n407), .C(buffer[253]), .D(n458), .Y(
        n987) );
  INVX1 U1241 ( .A(parallel_in[254]), .Y(n986) );
  OAI21X1 U1242 ( .A(n380), .B(n988), .C(n989), .Y(n1189) );
  AOI22X1 U1243 ( .A(buffer[255]), .B(n407), .C(buffer[254]), .D(n458), .Y(
        n989) );
  INVX1 U1244 ( .A(parallel_in[255]), .Y(n988) );
  OAI21X1 U1245 ( .A(n380), .B(n990), .C(n991), .Y(n1188) );
  AOI22X1 U1246 ( .A(buffer[256]), .B(n406), .C(buffer[255]), .D(n458), .Y(
        n991) );
  INVX1 U1247 ( .A(parallel_in[256]), .Y(n990) );
  OAI21X1 U1248 ( .A(n380), .B(n992), .C(n993), .Y(n1187) );
  AOI22X1 U1249 ( .A(buffer[257]), .B(n406), .C(buffer[256]), .D(n458), .Y(
        n993) );
  INVX1 U1250 ( .A(parallel_in[257]), .Y(n992) );
  OAI21X1 U1251 ( .A(n380), .B(n994), .C(n995), .Y(n1186) );
  AOI22X1 U1252 ( .A(buffer[258]), .B(n406), .C(buffer[257]), .D(n458), .Y(
        n995) );
  INVX1 U1253 ( .A(parallel_in[258]), .Y(n994) );
  OAI21X1 U1254 ( .A(n380), .B(n996), .C(n997), .Y(n1185) );
  AOI22X1 U1255 ( .A(buffer[259]), .B(n406), .C(buffer[258]), .D(n458), .Y(
        n997) );
  INVX1 U1256 ( .A(parallel_in[259]), .Y(n996) );
  OAI21X1 U1257 ( .A(n381), .B(n998), .C(n999), .Y(n1184) );
  AOI22X1 U1258 ( .A(buffer[260]), .B(n406), .C(buffer[259]), .D(n458), .Y(
        n999) );
  INVX1 U1259 ( .A(parallel_in[260]), .Y(n998) );
  OAI21X1 U1260 ( .A(n381), .B(n1000), .C(n1001), .Y(n1183) );
  AOI22X1 U1261 ( .A(buffer[261]), .B(n406), .C(buffer[260]), .D(n458), .Y(
        n1001) );
  INVX1 U1262 ( .A(parallel_in[261]), .Y(n1000) );
  OAI21X1 U1263 ( .A(n381), .B(n1002), .C(n1003), .Y(n1182) );
  AOI22X1 U1264 ( .A(buffer[262]), .B(n406), .C(buffer[261]), .D(n458), .Y(
        n1003) );
  INVX1 U1265 ( .A(parallel_in[262]), .Y(n1002) );
  OAI21X1 U1266 ( .A(n381), .B(n1004), .C(n1005), .Y(n1181) );
  AOI22X1 U1267 ( .A(buffer[263]), .B(n406), .C(buffer[262]), .D(n458), .Y(
        n1005) );
  INVX1 U1268 ( .A(parallel_in[263]), .Y(n1004) );
  OAI21X1 U1269 ( .A(n381), .B(n1006), .C(n1007), .Y(n1180) );
  AOI22X1 U1270 ( .A(buffer[264]), .B(n406), .C(buffer[263]), .D(n458), .Y(
        n1007) );
  INVX1 U1271 ( .A(parallel_in[264]), .Y(n1006) );
  OAI21X1 U1272 ( .A(n381), .B(n1008), .C(n1009), .Y(n1179) );
  AOI22X1 U1273 ( .A(buffer[265]), .B(n406), .C(buffer[264]), .D(n458), .Y(
        n1009) );
  INVX1 U1274 ( .A(parallel_in[265]), .Y(n1008) );
  OAI21X1 U1275 ( .A(n381), .B(n1010), .C(n1011), .Y(n1178) );
  AOI22X1 U1276 ( .A(buffer[266]), .B(n406), .C(buffer[265]), .D(n457), .Y(
        n1011) );
  INVX1 U1277 ( .A(parallel_in[266]), .Y(n1010) );
  OAI21X1 U1278 ( .A(n381), .B(n1012), .C(n1013), .Y(n1177) );
  AOI22X1 U1279 ( .A(buffer[267]), .B(n406), .C(buffer[266]), .D(n457), .Y(
        n1013) );
  INVX1 U1280 ( .A(parallel_in[267]), .Y(n1012) );
  OAI21X1 U1281 ( .A(n381), .B(n1014), .C(n1015), .Y(n1176) );
  AOI22X1 U1282 ( .A(buffer[268]), .B(n406), .C(buffer[267]), .D(n457), .Y(
        n1015) );
  INVX1 U1283 ( .A(parallel_in[268]), .Y(n1014) );
  OAI21X1 U1284 ( .A(n381), .B(n1016), .C(n1017), .Y(n1175) );
  AOI22X1 U1285 ( .A(buffer[269]), .B(n405), .C(buffer[268]), .D(n457), .Y(
        n1017) );
  INVX1 U1286 ( .A(parallel_in[269]), .Y(n1016) );
  OAI21X1 U1287 ( .A(n381), .B(n1018), .C(n1019), .Y(n1174) );
  AOI22X1 U1288 ( .A(buffer[270]), .B(n405), .C(buffer[269]), .D(n457), .Y(
        n1019) );
  INVX1 U1289 ( .A(parallel_in[270]), .Y(n1018) );
  OAI21X1 U1290 ( .A(n381), .B(n1020), .C(n1021), .Y(n1173) );
  AOI22X1 U1291 ( .A(buffer[271]), .B(n405), .C(buffer[270]), .D(n457), .Y(
        n1021) );
  INVX1 U1292 ( .A(parallel_in[271]), .Y(n1020) );
  OAI21X1 U1293 ( .A(n381), .B(n1022), .C(n1023), .Y(n1172) );
  AOI22X1 U1294 ( .A(buffer[272]), .B(n405), .C(buffer[271]), .D(n457), .Y(
        n1023) );
  INVX1 U1295 ( .A(parallel_in[272]), .Y(n1022) );
  OAI21X1 U1296 ( .A(n382), .B(n1024), .C(n1025), .Y(n1171) );
  AOI22X1 U1297 ( .A(buffer[273]), .B(n405), .C(buffer[272]), .D(n457), .Y(
        n1025) );
  INVX1 U1298 ( .A(parallel_in[273]), .Y(n1024) );
  OAI21X1 U1299 ( .A(n382), .B(n1026), .C(n1027), .Y(n1170) );
  AOI22X1 U1300 ( .A(buffer[274]), .B(n405), .C(buffer[273]), .D(n457), .Y(
        n1027) );
  INVX1 U1301 ( .A(parallel_in[274]), .Y(n1026) );
  OAI21X1 U1302 ( .A(n382), .B(n1028), .C(n1029), .Y(n1169) );
  AOI22X1 U1303 ( .A(buffer[275]), .B(n405), .C(buffer[274]), .D(n457), .Y(
        n1029) );
  INVX1 U1304 ( .A(parallel_in[275]), .Y(n1028) );
  OAI21X1 U1305 ( .A(n382), .B(n1030), .C(n1031), .Y(n1168) );
  AOI22X1 U1306 ( .A(buffer[276]), .B(n405), .C(buffer[275]), .D(n457), .Y(
        n1031) );
  INVX1 U1307 ( .A(parallel_in[276]), .Y(n1030) );
  OAI21X1 U1308 ( .A(n382), .B(n1032), .C(n1033), .Y(n1167) );
  AOI22X1 U1309 ( .A(buffer[277]), .B(n405), .C(buffer[276]), .D(n457), .Y(
        n1033) );
  INVX1 U1310 ( .A(parallel_in[277]), .Y(n1032) );
  OAI21X1 U1311 ( .A(n382), .B(n1034), .C(n1035), .Y(n1166) );
  AOI22X1 U1312 ( .A(buffer[278]), .B(n405), .C(buffer[277]), .D(n456), .Y(
        n1035) );
  INVX1 U1313 ( .A(parallel_in[278]), .Y(n1034) );
  OAI21X1 U1314 ( .A(n382), .B(n1036), .C(n1037), .Y(n1165) );
  AOI22X1 U1315 ( .A(buffer[279]), .B(n405), .C(buffer[278]), .D(n456), .Y(
        n1037) );
  INVX1 U1316 ( .A(parallel_in[279]), .Y(n1036) );
  OAI21X1 U1317 ( .A(n382), .B(n1038), .C(n1039), .Y(n1164) );
  AOI22X1 U1318 ( .A(buffer[280]), .B(n405), .C(buffer[279]), .D(n456), .Y(
        n1039) );
  INVX1 U1319 ( .A(parallel_in[280]), .Y(n1038) );
  OAI21X1 U1320 ( .A(n382), .B(n1040), .C(n1041), .Y(n1163) );
  AOI22X1 U1321 ( .A(buffer[281]), .B(n405), .C(buffer[280]), .D(n456), .Y(
        n1041) );
  INVX1 U1322 ( .A(parallel_in[281]), .Y(n1040) );
  OAI21X1 U1323 ( .A(n382), .B(n1042), .C(n1043), .Y(n1162) );
  AOI22X1 U1324 ( .A(buffer[282]), .B(n404), .C(buffer[281]), .D(n456), .Y(
        n1043) );
  INVX1 U1325 ( .A(parallel_in[282]), .Y(n1042) );
  OAI21X1 U1326 ( .A(n382), .B(n1044), .C(n1045), .Y(n1161) );
  AOI22X1 U1327 ( .A(buffer[283]), .B(n404), .C(buffer[282]), .D(n456), .Y(
        n1045) );
  INVX1 U1328 ( .A(parallel_in[283]), .Y(n1044) );
  OAI21X1 U1329 ( .A(n382), .B(n1046), .C(n1047), .Y(n1160) );
  AOI22X1 U1330 ( .A(buffer[284]), .B(n404), .C(buffer[283]), .D(n456), .Y(
        n1047) );
  INVX1 U1331 ( .A(parallel_in[284]), .Y(n1046) );
  OAI21X1 U1332 ( .A(n382), .B(n1048), .C(n1049), .Y(n1159) );
  AOI22X1 U1333 ( .A(buffer[285]), .B(n404), .C(buffer[284]), .D(n456), .Y(
        n1049) );
  INVX1 U1334 ( .A(parallel_in[285]), .Y(n1048) );
  OAI21X1 U1335 ( .A(n383), .B(n1050), .C(n1051), .Y(n1158) );
  AOI22X1 U1336 ( .A(buffer[286]), .B(n404), .C(buffer[285]), .D(n456), .Y(
        n1051) );
  INVX1 U1337 ( .A(parallel_in[286]), .Y(n1050) );
  OAI21X1 U1338 ( .A(n383), .B(n1052), .C(n1053), .Y(n1157) );
  AOI22X1 U1339 ( .A(buffer[287]), .B(n404), .C(buffer[286]), .D(n456), .Y(
        n1053) );
  INVX1 U1340 ( .A(parallel_in[287]), .Y(n1052) );
  OAI21X1 U1341 ( .A(n383), .B(n1054), .C(n1055), .Y(n1156) );
  AOI22X1 U1342 ( .A(buffer[288]), .B(n404), .C(buffer[287]), .D(n456), .Y(
        n1055) );
  INVX1 U1343 ( .A(parallel_in[288]), .Y(n1054) );
  OAI21X1 U1344 ( .A(n383), .B(n1056), .C(n1057), .Y(n1155) );
  AOI22X1 U1345 ( .A(buffer[289]), .B(n404), .C(buffer[288]), .D(n456), .Y(
        n1057) );
  INVX1 U1346 ( .A(parallel_in[289]), .Y(n1056) );
  OAI21X1 U1347 ( .A(n383), .B(n1058), .C(n1059), .Y(n1154) );
  AOI22X1 U1348 ( .A(buffer[290]), .B(n404), .C(buffer[289]), .D(n456), .Y(
        n1059) );
  INVX1 U1349 ( .A(parallel_in[290]), .Y(n1058) );
  OAI21X1 U1350 ( .A(n383), .B(n1060), .C(n1061), .Y(n1153) );
  AOI22X1 U1351 ( .A(buffer[291]), .B(n404), .C(buffer[290]), .D(n455), .Y(
        n1061) );
  INVX1 U1352 ( .A(parallel_in[291]), .Y(n1060) );
  OAI21X1 U1353 ( .A(n383), .B(n1062), .C(n1063), .Y(n1152) );
  AOI22X1 U1354 ( .A(buffer[292]), .B(n404), .C(buffer[291]), .D(n455), .Y(
        n1063) );
  INVX1 U1355 ( .A(parallel_in[292]), .Y(n1062) );
  OAI21X1 U1356 ( .A(n383), .B(n1064), .C(n1065), .Y(n1151) );
  AOI22X1 U1357 ( .A(buffer[293]), .B(n404), .C(buffer[292]), .D(n455), .Y(
        n1065) );
  INVX1 U1358 ( .A(parallel_in[293]), .Y(n1064) );
  OAI21X1 U1359 ( .A(n383), .B(n1066), .C(n1067), .Y(n1150) );
  AOI22X1 U1360 ( .A(buffer[294]), .B(n404), .C(buffer[293]), .D(n455), .Y(
        n1067) );
  INVX1 U1361 ( .A(parallel_in[294]), .Y(n1066) );
  OAI21X1 U1362 ( .A(n383), .B(n1068), .C(n1069), .Y(n1149) );
  AOI22X1 U1363 ( .A(buffer[295]), .B(n403), .C(buffer[294]), .D(n455), .Y(
        n1069) );
  INVX1 U1364 ( .A(parallel_in[295]), .Y(n1068) );
  OAI21X1 U1365 ( .A(n383), .B(n1070), .C(n1071), .Y(n1148) );
  AOI22X1 U1366 ( .A(buffer[296]), .B(n403), .C(buffer[295]), .D(n455), .Y(
        n1071) );
  INVX1 U1367 ( .A(parallel_in[296]), .Y(n1070) );
  OAI21X1 U1368 ( .A(n383), .B(n1072), .C(n1073), .Y(n1147) );
  AOI22X1 U1369 ( .A(buffer[297]), .B(n403), .C(buffer[296]), .D(n455), .Y(
        n1073) );
  INVX1 U1370 ( .A(parallel_in[297]), .Y(n1072) );
  OAI21X1 U1371 ( .A(n383), .B(n1074), .C(n1075), .Y(n1146) );
  AOI22X1 U1372 ( .A(buffer[298]), .B(n403), .C(buffer[297]), .D(n455), .Y(
        n1075) );
  INVX1 U1373 ( .A(parallel_in[298]), .Y(n1074) );
  OAI21X1 U1374 ( .A(n384), .B(n1076), .C(n1077), .Y(n1145) );
  AOI22X1 U1375 ( .A(buffer[299]), .B(n403), .C(buffer[298]), .D(n455), .Y(
        n1077) );
  INVX1 U1376 ( .A(parallel_in[299]), .Y(n1076) );
  OAI21X1 U1377 ( .A(n384), .B(n1078), .C(n1079), .Y(n1144) );
  AOI22X1 U1378 ( .A(buffer[300]), .B(n403), .C(buffer[299]), .D(n455), .Y(
        n1079) );
  INVX1 U1379 ( .A(parallel_in[300]), .Y(n1078) );
  OAI21X1 U1380 ( .A(n384), .B(n1080), .C(n1081), .Y(n1143) );
  AOI22X1 U1381 ( .A(buffer[301]), .B(n403), .C(buffer[300]), .D(n455), .Y(
        n1081) );
  INVX1 U1382 ( .A(parallel_in[301]), .Y(n1080) );
  OAI21X1 U1383 ( .A(n384), .B(n1082), .C(n1083), .Y(n1142) );
  AOI22X1 U1384 ( .A(buffer[302]), .B(n403), .C(buffer[301]), .D(n455), .Y(
        n1083) );
  INVX1 U1385 ( .A(parallel_in[302]), .Y(n1082) );
  OAI21X1 U1386 ( .A(n384), .B(n1084), .C(n1445), .Y(n1141) );
  AOI22X1 U1387 ( .A(buffer[303]), .B(n403), .C(buffer[302]), .D(n455), .Y(
        n1445) );
  INVX1 U1388 ( .A(parallel_in[303]), .Y(n1084) );
  OAI21X1 U1389 ( .A(n384), .B(n1446), .C(n1447), .Y(n1140) );
  AOI22X1 U1390 ( .A(buffer[304]), .B(n403), .C(buffer[303]), .D(n454), .Y(
        n1447) );
  INVX1 U1391 ( .A(parallel_in[304]), .Y(n1446) );
  OAI21X1 U1392 ( .A(n384), .B(n1448), .C(n1449), .Y(n1139) );
  AOI22X1 U1393 ( .A(buffer[305]), .B(n403), .C(buffer[304]), .D(n454), .Y(
        n1449) );
  INVX1 U1394 ( .A(parallel_in[305]), .Y(n1448) );
  OAI21X1 U1395 ( .A(n384), .B(n1450), .C(n1451), .Y(n1138) );
  AOI22X1 U1396 ( .A(buffer[306]), .B(n403), .C(buffer[305]), .D(n454), .Y(
        n1451) );
  INVX1 U1397 ( .A(parallel_in[306]), .Y(n1450) );
  OAI21X1 U1398 ( .A(n384), .B(n1452), .C(n1453), .Y(n1137) );
  AOI22X1 U1399 ( .A(buffer[307]), .B(n403), .C(buffer[306]), .D(n454), .Y(
        n1453) );
  INVX1 U1400 ( .A(parallel_in[307]), .Y(n1452) );
  OAI21X1 U1401 ( .A(n384), .B(n1454), .C(n1455), .Y(n1136) );
  AOI22X1 U1402 ( .A(buffer[308]), .B(n402), .C(buffer[307]), .D(n454), .Y(
        n1455) );
  INVX1 U1403 ( .A(parallel_in[308]), .Y(n1454) );
  OAI21X1 U1404 ( .A(n384), .B(n1456), .C(n1457), .Y(n1135) );
  AOI22X1 U1405 ( .A(buffer[309]), .B(n402), .C(buffer[308]), .D(n454), .Y(
        n1457) );
  INVX1 U1406 ( .A(parallel_in[309]), .Y(n1456) );
  OAI21X1 U1407 ( .A(n384), .B(n1458), .C(n1459), .Y(n1134) );
  AOI22X1 U1408 ( .A(buffer[310]), .B(n402), .C(buffer[309]), .D(n454), .Y(
        n1459) );
  INVX1 U1409 ( .A(parallel_in[310]), .Y(n1458) );
  OAI21X1 U1410 ( .A(n384), .B(n1460), .C(n1461), .Y(n1133) );
  AOI22X1 U1411 ( .A(buffer[311]), .B(n402), .C(buffer[310]), .D(n454), .Y(
        n1461) );
  INVX1 U1412 ( .A(parallel_in[311]), .Y(n1460) );
  OAI21X1 U1413 ( .A(n385), .B(n1462), .C(n1463), .Y(n1132) );
  AOI22X1 U1414 ( .A(buffer[312]), .B(n402), .C(buffer[311]), .D(n454), .Y(
        n1463) );
  INVX1 U1415 ( .A(parallel_in[312]), .Y(n1462) );
  OAI21X1 U1416 ( .A(n385), .B(n1464), .C(n1465), .Y(n1131) );
  AOI22X1 U1417 ( .A(buffer[313]), .B(n402), .C(buffer[312]), .D(n454), .Y(
        n1465) );
  INVX1 U1418 ( .A(parallel_in[313]), .Y(n1464) );
  OAI21X1 U1419 ( .A(n385), .B(n1466), .C(n1467), .Y(n1130) );
  AOI22X1 U1420 ( .A(buffer[314]), .B(n402), .C(buffer[313]), .D(n454), .Y(
        n1467) );
  INVX1 U1421 ( .A(parallel_in[314]), .Y(n1466) );
  OAI21X1 U1422 ( .A(n385), .B(n1468), .C(n1469), .Y(n1129) );
  AOI22X1 U1423 ( .A(buffer[315]), .B(n402), .C(buffer[314]), .D(n454), .Y(
        n1469) );
  INVX1 U1424 ( .A(parallel_in[315]), .Y(n1468) );
  OAI21X1 U1425 ( .A(n385), .B(n1470), .C(n1471), .Y(n1128) );
  AOI22X1 U1426 ( .A(buffer[316]), .B(n402), .C(buffer[315]), .D(n454), .Y(
        n1471) );
  INVX1 U1427 ( .A(parallel_in[316]), .Y(n1470) );
  OAI21X1 U1428 ( .A(n385), .B(n1472), .C(n1473), .Y(n1127) );
  AOI22X1 U1429 ( .A(buffer[317]), .B(n402), .C(buffer[316]), .D(n453), .Y(
        n1473) );
  INVX1 U1430 ( .A(parallel_in[317]), .Y(n1472) );
  OAI21X1 U1431 ( .A(n385), .B(n1474), .C(n1475), .Y(n1126) );
  AOI22X1 U1432 ( .A(buffer[318]), .B(n402), .C(buffer[317]), .D(n457), .Y(
        n1475) );
  INVX1 U1433 ( .A(parallel_in[318]), .Y(n1474) );
  OAI21X1 U1434 ( .A(n385), .B(n1476), .C(n1477), .Y(n1125) );
  AOI22X1 U1435 ( .A(buffer[319]), .B(n402), .C(buffer[318]), .D(n453), .Y(
        n1477) );
  INVX1 U1436 ( .A(parallel_in[319]), .Y(n1476) );
  OAI21X1 U1437 ( .A(n385), .B(n1478), .C(n1479), .Y(n1124) );
  AOI22X1 U1438 ( .A(buffer[320]), .B(n402), .C(buffer[319]), .D(n453), .Y(
        n1479) );
  INVX1 U1439 ( .A(parallel_in[320]), .Y(n1478) );
  OAI21X1 U1440 ( .A(n385), .B(n1480), .C(n1481), .Y(n1123) );
  AOI22X1 U1441 ( .A(buffer[321]), .B(n401), .C(buffer[320]), .D(n453), .Y(
        n1481) );
  INVX1 U1442 ( .A(parallel_in[321]), .Y(n1480) );
  OAI21X1 U1443 ( .A(n385), .B(n1482), .C(n1483), .Y(n1122) );
  AOI22X1 U1444 ( .A(buffer[322]), .B(n401), .C(buffer[321]), .D(n453), .Y(
        n1483) );
  INVX1 U1445 ( .A(parallel_in[322]), .Y(n1482) );
  OAI21X1 U1446 ( .A(n385), .B(n1484), .C(n1485), .Y(n1121) );
  AOI22X1 U1447 ( .A(buffer[323]), .B(n401), .C(buffer[322]), .D(n453), .Y(
        n1485) );
  INVX1 U1448 ( .A(parallel_in[323]), .Y(n1484) );
  OAI21X1 U1449 ( .A(n385), .B(n1486), .C(n1487), .Y(n1120) );
  AOI22X1 U1450 ( .A(buffer[324]), .B(n401), .C(buffer[323]), .D(n453), .Y(
        n1487) );
  INVX1 U1451 ( .A(parallel_in[324]), .Y(n1486) );
  OAI21X1 U1452 ( .A(n386), .B(n1488), .C(n1489), .Y(n1119) );
  AOI22X1 U1453 ( .A(buffer[325]), .B(n401), .C(buffer[324]), .D(n453), .Y(
        n1489) );
  INVX1 U1454 ( .A(parallel_in[325]), .Y(n1488) );
  OAI21X1 U1455 ( .A(n386), .B(n1490), .C(n1491), .Y(n1118) );
  AOI22X1 U1456 ( .A(buffer[326]), .B(n401), .C(buffer[325]), .D(n453), .Y(
        n1491) );
  INVX1 U1457 ( .A(parallel_in[326]), .Y(n1490) );
  OAI21X1 U1458 ( .A(n386), .B(n1492), .C(n1493), .Y(n1117) );
  AOI22X1 U1459 ( .A(buffer[327]), .B(n401), .C(buffer[326]), .D(n453), .Y(
        n1493) );
  INVX1 U1460 ( .A(parallel_in[327]), .Y(n1492) );
  OAI21X1 U1461 ( .A(n386), .B(n1494), .C(n1495), .Y(n1116) );
  AOI22X1 U1462 ( .A(buffer[328]), .B(n401), .C(buffer[327]), .D(n453), .Y(
        n1495) );
  INVX1 U1463 ( .A(parallel_in[328]), .Y(n1494) );
  OAI21X1 U1464 ( .A(n386), .B(n1496), .C(n1497), .Y(n1115) );
  AOI22X1 U1465 ( .A(buffer[329]), .B(n401), .C(buffer[328]), .D(n453), .Y(
        n1497) );
  INVX1 U1466 ( .A(parallel_in[329]), .Y(n1496) );
  OAI21X1 U1467 ( .A(n386), .B(n1498), .C(n1499), .Y(n1114) );
  AOI22X1 U1468 ( .A(buffer[330]), .B(n401), .C(buffer[329]), .D(n453), .Y(
        n1499) );
  INVX1 U1469 ( .A(parallel_in[330]), .Y(n1498) );
  OAI21X1 U1470 ( .A(n386), .B(n1500), .C(n1501), .Y(n1113) );
  AOI22X1 U1471 ( .A(buffer[331]), .B(n401), .C(buffer[330]), .D(n452), .Y(
        n1501) );
  INVX1 U1472 ( .A(parallel_in[331]), .Y(n1500) );
  OAI21X1 U1473 ( .A(n386), .B(n1502), .C(n1503), .Y(n1112) );
  AOI22X1 U1474 ( .A(buffer[332]), .B(n401), .C(buffer[331]), .D(n452), .Y(
        n1503) );
  INVX1 U1475 ( .A(parallel_in[332]), .Y(n1502) );
  OAI21X1 U1476 ( .A(n386), .B(n1504), .C(n1505), .Y(n1111) );
  AOI22X1 U1477 ( .A(buffer[333]), .B(n401), .C(buffer[332]), .D(n452), .Y(
        n1505) );
  INVX1 U1478 ( .A(parallel_in[333]), .Y(n1504) );
  OAI21X1 U1479 ( .A(n386), .B(n1506), .C(n1507), .Y(n1110) );
  AOI22X1 U1480 ( .A(buffer[334]), .B(n400), .C(buffer[333]), .D(n452), .Y(
        n1507) );
  INVX1 U1481 ( .A(parallel_in[334]), .Y(n1506) );
  OAI21X1 U1482 ( .A(n386), .B(n1508), .C(n1509), .Y(n1109) );
  AOI22X1 U1483 ( .A(buffer[335]), .B(n400), .C(buffer[334]), .D(n452), .Y(
        n1509) );
  INVX1 U1484 ( .A(parallel_in[335]), .Y(n1508) );
  OAI21X1 U1485 ( .A(n386), .B(n1510), .C(n1511), .Y(n1108) );
  AOI22X1 U1486 ( .A(buffer[336]), .B(n400), .C(buffer[335]), .D(n452), .Y(
        n1511) );
  INVX1 U1487 ( .A(parallel_in[336]), .Y(n1510) );
  OAI21X1 U1488 ( .A(n386), .B(n1512), .C(n1513), .Y(n1107) );
  AOI22X1 U1489 ( .A(buffer[337]), .B(n400), .C(buffer[336]), .D(n452), .Y(
        n1513) );
  INVX1 U1490 ( .A(parallel_in[337]), .Y(n1512) );
  OAI21X1 U1491 ( .A(n387), .B(n1514), .C(n1515), .Y(n1106) );
  AOI22X1 U1492 ( .A(buffer[338]), .B(n400), .C(buffer[337]), .D(n452), .Y(
        n1515) );
  INVX1 U1493 ( .A(parallel_in[338]), .Y(n1514) );
  OAI21X1 U1494 ( .A(n387), .B(n1516), .C(n1517), .Y(n1105) );
  AOI22X1 U1495 ( .A(buffer[339]), .B(n400), .C(buffer[338]), .D(n452), .Y(
        n1517) );
  INVX1 U1496 ( .A(parallel_in[339]), .Y(n1516) );
  OAI21X1 U1497 ( .A(n387), .B(n1518), .C(n1519), .Y(n1104) );
  AOI22X1 U1498 ( .A(buffer[340]), .B(n400), .C(buffer[339]), .D(n452), .Y(
        n1519) );
  INVX1 U1499 ( .A(parallel_in[340]), .Y(n1518) );
  OAI21X1 U1500 ( .A(n387), .B(n1520), .C(n1521), .Y(n1103) );
  AOI22X1 U1501 ( .A(buffer[341]), .B(n400), .C(buffer[340]), .D(n452), .Y(
        n1521) );
  INVX1 U1502 ( .A(parallel_in[341]), .Y(n1520) );
  OAI21X1 U1503 ( .A(n387), .B(n1522), .C(n1523), .Y(n1102) );
  AOI22X1 U1504 ( .A(buffer[342]), .B(n400), .C(buffer[341]), .D(n452), .Y(
        n1523) );
  INVX1 U1505 ( .A(parallel_in[342]), .Y(n1522) );
  OAI21X1 U1506 ( .A(n387), .B(n1524), .C(n1525), .Y(n1101) );
  AOI22X1 U1507 ( .A(buffer[343]), .B(n400), .C(buffer[342]), .D(n452), .Y(
        n1525) );
  INVX1 U1508 ( .A(parallel_in[343]), .Y(n1524) );
  OAI21X1 U1509 ( .A(n387), .B(n1526), .C(n1527), .Y(n1100) );
  AOI22X1 U1510 ( .A(buffer[344]), .B(n400), .C(buffer[343]), .D(n451), .Y(
        n1527) );
  INVX1 U1511 ( .A(parallel_in[344]), .Y(n1526) );
  OAI21X1 U1512 ( .A(n387), .B(n1528), .C(n1529), .Y(n1099) );
  AOI22X1 U1513 ( .A(buffer[345]), .B(n400), .C(buffer[344]), .D(n451), .Y(
        n1529) );
  INVX1 U1514 ( .A(parallel_in[345]), .Y(n1528) );
  OAI21X1 U1515 ( .A(n387), .B(n1530), .C(n1531), .Y(n1098) );
  AOI22X1 U1516 ( .A(buffer[346]), .B(n400), .C(buffer[345]), .D(n451), .Y(
        n1531) );
  INVX1 U1517 ( .A(parallel_in[346]), .Y(n1530) );
  OAI21X1 U1518 ( .A(n387), .B(n1532), .C(n1533), .Y(n1097) );
  AOI22X1 U1519 ( .A(buffer[347]), .B(n399), .C(buffer[346]), .D(n451), .Y(
        n1533) );
  INVX1 U1520 ( .A(parallel_in[347]), .Y(n1532) );
  OAI21X1 U1521 ( .A(n387), .B(n1534), .C(n1535), .Y(n1096) );
  AOI22X1 U1522 ( .A(buffer[348]), .B(n399), .C(buffer[347]), .D(n451), .Y(
        n1535) );
  INVX1 U1523 ( .A(parallel_in[348]), .Y(n1534) );
  OAI21X1 U1524 ( .A(n387), .B(n1536), .C(n1537), .Y(n1095) );
  AOI22X1 U1525 ( .A(buffer[349]), .B(n399), .C(buffer[348]), .D(n451), .Y(
        n1537) );
  INVX1 U1526 ( .A(parallel_in[349]), .Y(n1536) );
  OAI21X1 U1527 ( .A(n387), .B(n1538), .C(n1539), .Y(n1094) );
  AOI22X1 U1528 ( .A(buffer[350]), .B(n399), .C(buffer[349]), .D(n451), .Y(
        n1539) );
  INVX1 U1529 ( .A(parallel_in[350]), .Y(n1538) );
  OAI21X1 U1530 ( .A(n388), .B(n1540), .C(n1541), .Y(n1093) );
  AOI22X1 U1531 ( .A(buffer[351]), .B(n399), .C(buffer[350]), .D(n451), .Y(
        n1541) );
  INVX1 U1532 ( .A(parallel_in[351]), .Y(n1540) );
  OAI21X1 U1533 ( .A(n388), .B(n1542), .C(n1543), .Y(n1092) );
  AOI22X1 U1534 ( .A(buffer[352]), .B(n399), .C(buffer[351]), .D(n451), .Y(
        n1543) );
  INVX1 U1535 ( .A(parallel_in[352]), .Y(n1542) );
  OAI21X1 U1536 ( .A(n388), .B(n1544), .C(n1545), .Y(n1091) );
  AOI22X1 U1537 ( .A(buffer[353]), .B(n399), .C(buffer[352]), .D(n451), .Y(
        n1545) );
  INVX1 U1538 ( .A(parallel_in[353]), .Y(n1544) );
  OAI21X1 U1539 ( .A(n388), .B(n1546), .C(n1547), .Y(n1090) );
  AOI22X1 U1540 ( .A(buffer[354]), .B(n399), .C(buffer[353]), .D(n451), .Y(
        n1547) );
  INVX1 U1541 ( .A(parallel_in[354]), .Y(n1546) );
  OAI21X1 U1542 ( .A(n388), .B(n1548), .C(n1549), .Y(n1089) );
  AOI22X1 U1543 ( .A(buffer[355]), .B(n399), .C(buffer[354]), .D(n451), .Y(
        n1549) );
  INVX1 U1544 ( .A(parallel_in[355]), .Y(n1548) );
  OAI21X1 U1545 ( .A(n388), .B(n1550), .C(n1551), .Y(n1088) );
  AOI22X1 U1546 ( .A(buffer[356]), .B(n399), .C(buffer[355]), .D(n451), .Y(
        n1551) );
  INVX1 U1547 ( .A(parallel_in[356]), .Y(n1550) );
  OAI21X1 U1548 ( .A(n388), .B(n1552), .C(n1553), .Y(n1087) );
  AOI22X1 U1549 ( .A(buffer[357]), .B(n399), .C(buffer[356]), .D(n450), .Y(
        n1553) );
  INVX1 U1550 ( .A(parallel_in[357]), .Y(n1552) );
  OAI21X1 U1551 ( .A(n388), .B(n1554), .C(n1555), .Y(n1086) );
  AOI22X1 U1552 ( .A(buffer[358]), .B(n399), .C(buffer[357]), .D(n450), .Y(
        n1555) );
  INVX1 U1553 ( .A(parallel_in[358]), .Y(n1554) );
  OAI21X1 U1554 ( .A(n388), .B(n1556), .C(n1557), .Y(n1085) );
  AOI22X1 U1555 ( .A(serial_out), .B(n399), .C(buffer[358]), .D(n450), .Y(
        n1557) );
  NOR2X1 U1556 ( .A(load_enable), .B(n464), .Y(n478) );
  AND2X1 U1557 ( .A(shift_enable), .B(n388), .Y(n479) );
  INVX1 U1558 ( .A(parallel_in[359]), .Y(n1556) );
  INVX1 U1559 ( .A(load_enable), .Y(n476) );
endmodule


module flex_counter_NUM_CNT_BITS9_DW01_inc_0 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HAX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  HAX1 U1_1_6 ( .A(A[6]), .B(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  HAX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .YC(carry[6]), .YS(SUM[5]) );
  HAX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .YC(carry[5]), .YS(SUM[4]) );
  HAX1 U1_1_3 ( .A(A[3]), .B(carry[3]), .YC(carry[4]), .YS(SUM[3]) );
  HAX1 U1_1_2 ( .A(A[2]), .B(carry[2]), .YC(carry[3]), .YS(SUM[2]) );
  HAX1 U1_1_1 ( .A(A[1]), .B(A[0]), .YC(carry[2]), .YS(SUM[1]) );
  INVX2 U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1 U2 ( .A(carry[8]), .B(A[8]), .Y(SUM[8]) );
endmodule


module flex_counter_NUM_CNT_BITS9 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [8:0] rollover_val;
  output [8:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N22, \eq_50/A[0] ,
         \eq_50/A[1] , \eq_50/A[2] , \eq_50/A[3] , \eq_50/A[4] , \eq_50/A[5] ,
         \eq_50/A[6] , \eq_50/A[7] , \eq_50/A[8] , n1, n2, n3, n4, n5, n6, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62;

  DFFSR \count_out_reg[0]  ( .D(\eq_50/A[0] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[0]) );
  DFFSR \count_out_reg[8]  ( .D(\eq_50/A[8] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[8]) );
  DFFSR \count_out_reg[7]  ( .D(\eq_50/A[7] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[7]) );
  DFFSR \count_out_reg[6]  ( .D(\eq_50/A[6] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[6]) );
  DFFSR \count_out_reg[5]  ( .D(\eq_50/A[5] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[5]) );
  DFFSR \count_out_reg[4]  ( .D(\eq_50/A[4] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[4]) );
  DFFSR \count_out_reg[3]  ( .D(\eq_50/A[3] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[3]) );
  DFFSR \count_out_reg[2]  ( .D(\eq_50/A[2] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[2]) );
  DFFSR \count_out_reg[1]  ( .D(\eq_50/A[1] ), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[1]) );
  DFFSR rollover_flag_reg ( .D(N22), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        rollover_flag) );
  flex_counter_NUM_CNT_BITS9_DW01_inc_0 add_46 ( .A(count_out), .SUM({N15, N14, 
        N13, N12, N11, N10, N9, N8, N7}) );
  NOR2X1 U5 ( .A(n1), .B(n2), .Y(N22) );
  NAND3X1 U6 ( .A(n3), .B(n4), .C(n5), .Y(n2) );
  NOR2X1 U15 ( .A(n6), .B(n17), .Y(n5) );
  XOR2X1 U16 ( .A(rollover_val[8]), .B(\eq_50/A[8] ), .Y(n6) );
  OAI21X1 U17 ( .A(n18), .B(n19), .C(n20), .Y(\eq_50/A[8] ) );
  NAND2X1 U18 ( .A(N15), .B(n21), .Y(n20) );
  XNOR2X1 U19 ( .A(rollover_val[7]), .B(\eq_50/A[7] ), .Y(n4) );
  OAI21X1 U20 ( .A(n22), .B(n19), .C(n23), .Y(\eq_50/A[7] ) );
  NAND2X1 U21 ( .A(N14), .B(n21), .Y(n23) );
  NOR2X1 U22 ( .A(n24), .B(n25), .Y(n3) );
  XOR2X1 U23 ( .A(rollover_val[4]), .B(\eq_50/A[4] ), .Y(n25) );
  OAI21X1 U24 ( .A(n26), .B(n19), .C(n27), .Y(\eq_50/A[4] ) );
  NAND2X1 U25 ( .A(N11), .B(n21), .Y(n27) );
  INVX1 U26 ( .A(count_out[4]), .Y(n26) );
  XOR2X1 U27 ( .A(rollover_val[5]), .B(\eq_50/A[5] ), .Y(n24) );
  OAI21X1 U28 ( .A(n28), .B(n19), .C(n29), .Y(\eq_50/A[5] ) );
  NAND2X1 U29 ( .A(N12), .B(n21), .Y(n29) );
  INVX1 U30 ( .A(count_out[5]), .Y(n28) );
  NAND3X1 U31 ( .A(n30), .B(n31), .C(n32), .Y(n1) );
  NOR2X1 U32 ( .A(n33), .B(n34), .Y(n32) );
  XOR2X1 U33 ( .A(rollover_val[6]), .B(\eq_50/A[6] ), .Y(n34) );
  OAI21X1 U34 ( .A(n35), .B(n19), .C(n36), .Y(\eq_50/A[6] ) );
  NAND2X1 U35 ( .A(N13), .B(n21), .Y(n36) );
  INVX1 U36 ( .A(count_out[6]), .Y(n35) );
  XOR2X1 U37 ( .A(rollover_val[3]), .B(\eq_50/A[3] ), .Y(n33) );
  OAI21X1 U38 ( .A(n37), .B(n19), .C(n38), .Y(\eq_50/A[3] ) );
  NAND2X1 U39 ( .A(N10), .B(n21), .Y(n38) );
  INVX1 U40 ( .A(count_out[3]), .Y(n37) );
  XNOR2X1 U41 ( .A(rollover_val[2]), .B(\eq_50/A[2] ), .Y(n31) );
  OAI21X1 U42 ( .A(n39), .B(n19), .C(n40), .Y(\eq_50/A[2] ) );
  NAND2X1 U43 ( .A(N9), .B(n21), .Y(n40) );
  INVX1 U44 ( .A(count_out[2]), .Y(n39) );
  NOR2X1 U45 ( .A(n41), .B(n42), .Y(n30) );
  XOR2X1 U46 ( .A(rollover_val[0]), .B(\eq_50/A[0] ), .Y(n42) );
  OAI21X1 U47 ( .A(n43), .B(n19), .C(n44), .Y(\eq_50/A[0] ) );
  NAND2X1 U48 ( .A(N7), .B(n21), .Y(n44) );
  INVX1 U49 ( .A(count_out[0]), .Y(n43) );
  XOR2X1 U50 ( .A(rollover_val[1]), .B(\eq_50/A[1] ), .Y(n41) );
  OAI21X1 U51 ( .A(n45), .B(n19), .C(n46), .Y(\eq_50/A[1] ) );
  NAND2X1 U52 ( .A(N8), .B(n21), .Y(n46) );
  NOR2X1 U53 ( .A(n17), .B(n47), .Y(n21) );
  OAI21X1 U54 ( .A(n48), .B(n49), .C(n50), .Y(n47) );
  NAND3X1 U55 ( .A(n51), .B(n52), .C(n53), .Y(n49) );
  NOR2X1 U56 ( .A(n54), .B(n55), .Y(n53) );
  XOR2X1 U57 ( .A(rollover_val[6]), .B(count_out[6]), .Y(n55) );
  XOR2X1 U58 ( .A(rollover_val[5]), .B(count_out[5]), .Y(n54) );
  XOR2X1 U59 ( .A(n22), .B(rollover_val[7]), .Y(n52) );
  INVX1 U60 ( .A(count_out[7]), .Y(n22) );
  XOR2X1 U61 ( .A(n18), .B(rollover_val[8]), .Y(n51) );
  INVX1 U62 ( .A(count_out[8]), .Y(n18) );
  NAND3X1 U63 ( .A(n56), .B(n57), .C(n58), .Y(n48) );
  NOR2X1 U64 ( .A(n59), .B(n60), .Y(n58) );
  XOR2X1 U65 ( .A(rollover_val[4]), .B(count_out[4]), .Y(n60) );
  XOR2X1 U66 ( .A(rollover_val[3]), .B(count_out[3]), .Y(n59) );
  XOR2X1 U67 ( .A(n45), .B(rollover_val[1]), .Y(n57) );
  NOR2X1 U68 ( .A(n61), .B(n62), .Y(n56) );
  XOR2X1 U69 ( .A(rollover_val[0]), .B(count_out[0]), .Y(n62) );
  XOR2X1 U70 ( .A(rollover_val[2]), .B(count_out[2]), .Y(n61) );
  NAND2X1 U71 ( .A(n17), .B(n50), .Y(n19) );
  INVX1 U72 ( .A(clear), .Y(n50) );
  INVX1 U73 ( .A(count_enable), .Y(n17) );
  INVX1 U74 ( .A(count_out[1]), .Y(n45) );
endmodule


module flex_counter_NUM_CNT_BITS4 ( clk, n_rst, clear, count_enable, 
        rollover_val, count_out, rollover_flag );
  input [3:0] rollover_val;
  output [3:0] count_out;
  input clk, n_rst, clear, count_enable;
  output rollover_flag;
  wire   n1, n2, n3, n4, n5, n6, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35;
  wire   [3:0] nxt_data;

  DFFSR \count_out_reg[0]  ( .D(nxt_data[0]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[0]) );
  DFFSR \count_out_reg[1]  ( .D(nxt_data[1]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[1]) );
  DFFSR \count_out_reg[3]  ( .D(nxt_data[3]), .CLK(clk), .R(n_rst), .S(1'b1), 
        .Q(count_out[3]) );
  DFFSR \count_out_reg[2]  ( .D(n35), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        count_out[2]) );
  DFFSR rollover_flag_reg ( .D(n34), .CLK(clk), .R(n_rst), .S(1'b1), .Q(
        rollover_flag) );
  INVX1 U8 ( .A(n1), .Y(n34) );
  NAND3X1 U9 ( .A(n2), .B(n3), .C(n4), .Y(n1) );
  NOR2X1 U10 ( .A(n5), .B(n6), .Y(n4) );
  OAI21X1 U11 ( .A(nxt_data[0]), .B(n12), .C(n13), .Y(n6) );
  XNOR2X1 U12 ( .A(rollover_val[2]), .B(n35), .Y(n13) );
  MUX2X1 U13 ( .B(n14), .A(n15), .S(count_out[0]), .Y(nxt_data[0]) );
  NAND2X1 U14 ( .A(n5), .B(n16), .Y(n15) );
  XNOR2X1 U15 ( .A(nxt_data[1]), .B(rollover_val[1]), .Y(n3) );
  MUX2X1 U16 ( .B(n17), .A(n18), .S(count_out[1]), .Y(nxt_data[1]) );
  NAND2X1 U17 ( .A(count_out[0]), .B(n19), .Y(n17) );
  XNOR2X1 U18 ( .A(nxt_data[3]), .B(rollover_val[3]), .Y(n2) );
  INVX1 U19 ( .A(n20), .Y(nxt_data[3]) );
  MUX2X1 U20 ( .B(n21), .A(n22), .S(count_out[3]), .Y(n20) );
  OAI21X1 U21 ( .A(count_out[2]), .B(n14), .C(n23), .Y(n22) );
  NOR2X1 U22 ( .A(n24), .B(n25), .Y(n21) );
  MUX2X1 U23 ( .B(n23), .A(n25), .S(n24), .Y(n35) );
  INVX1 U24 ( .A(count_out[2]), .Y(n24) );
  NAND3X1 U25 ( .A(count_out[1]), .B(count_out[0]), .C(n19), .Y(n25) );
  INVX1 U26 ( .A(n26), .Y(n23) );
  OAI21X1 U27 ( .A(count_out[1]), .B(n14), .C(n18), .Y(n26) );
  AOI22X1 U28 ( .A(n5), .B(n16), .C(n27), .D(n19), .Y(n18) );
  INVX1 U29 ( .A(n14), .Y(n19) );
  INVX1 U30 ( .A(count_out[0]), .Y(n27) );
  INVX1 U31 ( .A(count_enable), .Y(n5) );
  NAND3X1 U32 ( .A(n28), .B(n16), .C(count_enable), .Y(n14) );
  INVX1 U33 ( .A(clear), .Y(n16) );
  NAND3X1 U34 ( .A(n29), .B(n30), .C(n31), .Y(n28) );
  NOR2X1 U35 ( .A(n32), .B(n33), .Y(n31) );
  XOR2X1 U36 ( .A(rollover_val[1]), .B(count_out[1]), .Y(n33) );
  XNOR2X1 U37 ( .A(n12), .B(count_out[0]), .Y(n32) );
  INVX1 U38 ( .A(rollover_val[0]), .Y(n12) );
  XNOR2X1 U39 ( .A(rollover_val[2]), .B(count_out[2]), .Y(n30) );
  XNOR2X1 U40 ( .A(count_out[3]), .B(rollover_val[3]), .Y(n29) );
endmodule


module uart_tx2 ( clk, n_rst, tx_data, send_data, serial_out );
  input [287:0] tx_data;
  input clk, n_rst, send_data;
  output serial_out;
  wire   done, tim_en, load_en, shift_enable;

  uart_tx_TCU UTT2 ( .clk(clk), .n_rst(n_rst), .send_data(send_data), .done(
        done), .tim_en(tim_en), .load_en(load_en) );
  flex_pts_sr_NUM_BITS360_SHIFT_MSB1 FPS2 ( .clk(clk), .n_rst(n_rst), 
        .shift_enable(shift_enable), .load_enable(load_en), .parallel_in({1'b0, 
        tx_data[287:280], 1'b1, 1'b0, tx_data[279:272], 1'b1, 1'b0, 
        tx_data[271:264], 1'b1, 1'b0, tx_data[263:256], 1'b1, 1'b0, 
        tx_data[255:248], 1'b1, 1'b0, tx_data[247:240], 1'b1, 1'b0, 
        tx_data[239:232], 1'b1, 1'b0, tx_data[231:224], 1'b1, 1'b0, 
        tx_data[223:216], 1'b1, 1'b0, tx_data[215:208], 1'b1, 1'b0, 
        tx_data[207:200], 1'b1, 1'b0, tx_data[199:192], 1'b1, 1'b0, 
        tx_data[191:184], 1'b1, 1'b0, tx_data[183:176], 1'b1, 1'b0, 
        tx_data[175:168], 1'b1, 1'b0, tx_data[167:160], 1'b1, 1'b0, 
        tx_data[159:152], 1'b1, 1'b0, tx_data[151:144], 1'b1, 1'b0, 
        tx_data[143:136], 1'b1, 1'b0, tx_data[135:128], 1'b1, 1'b0, 
        tx_data[127:120], 1'b1, 1'b0, tx_data[119:112], 1'b1, 1'b0, 
        tx_data[111:104], 1'b1, 1'b0, tx_data[103:96], 1'b1, 1'b0, 
        tx_data[95:88], 1'b1, 1'b0, tx_data[87:80], 1'b1, 1'b0, tx_data[79:72], 
        1'b1, 1'b0, tx_data[71:64], 1'b1, 1'b0, tx_data[63:56], 1'b1, 1'b0, 
        tx_data[55:48], 1'b1, 1'b0, tx_data[47:40], 1'b1, 1'b0, tx_data[39:32], 
        1'b1, 1'b0, tx_data[31:24], 1'b1, 1'b0, tx_data[23:16], 1'b1, 1'b0, 
        tx_data[15:8], 1'b1, 1'b0, tx_data[7:0], 1'b1}), .serial_out(
        serial_out) );
  flex_counter_NUM_CNT_BITS9 FC5 ( .clk(clk), .n_rst(n_rst), .clear(send_data), 
        .count_enable(shift_enable), .rollover_val({1'b1, 1'b0, 1'b1, 1'b1, 
        1'b0, 1'b1, 1'b0, 1'b0, 1'b0}), .rollover_flag(done) );
  flex_counter_NUM_CNT_BITS4 FC4 ( .clk(clk), .n_rst(n_rst), .clear(send_data), 
        .count_enable(tim_en), .rollover_val({1'b1, 1'b0, 1'b1, 1'b0}), 
        .rollover_flag(shift_enable) );
endmodule

