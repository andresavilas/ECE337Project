library verilog;
use verilog.vl_types.all;
entity tb_miner_core_comp is
end tb_miner_core_comp;
