library verilog;
use verilog.vl_types.all;
entity tb_bitcoinminer_sv_unit is
end tb_bitcoinminer_sv_unit;
