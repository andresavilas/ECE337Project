library verilog;
use verilog.vl_types.all;
entity tb_bitcoinminer is
end tb_bitcoinminer;
