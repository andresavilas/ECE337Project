library verilog;
use verilog.vl_types.all;
entity tb_miner is
end tb_miner;
