// $Id: $
// File name:   miner_core_msa.sv
// Created:     4/16/2015
// Author:      Andres Avila
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Message Scheduling Array
module miner_core_msa (
  input wire msa_en,
  input wire clk,
  input wire n_rst,
  input wire [0:511] chunk,
  output logic [0:63] [0:31] w 
);
  logic [0:31] s0;
  logic [0:31] s1;
  logic [0:31] w16;
  logic [0:31] w7;
  logic [0:31] w15;
  logic [0:31] w2;
  logic [0:31] out;
  logic [0:63] [0:31] new_w;
  reg [0:6] next_state;
  reg [0:6] state;
  always_ff @ (posedge clk, negedge n_rst) begin
    if(n_rst == 0) begin
      w <= 0;
      state <= 15;
    end else begin
      w <= new_w;
      state <= next_state;
    end
  end 
  always_comb begin
    next_state = state;
    new_w = w;
    case (state) 
  15: begin
    if(msa_en == 1) begin
      next_state = 16;
      new_w[0:15] = chunk;
    end 
  end
    16: begin
    w15 = w[1];
    w2 = w[14];
    w16 = w[0];
    w7 = w[9];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[16] = w16 + s0 + s1 + w7;
  end
  17: begin
    w15 = w[2];
    w2 = w[15];
    w16 = w[1];
    w7 = w[10];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[17] = w16 + s0 + s1 + w7;
  end
  18: begin
    w15 = w[3];
    w2 = w[16];
    w16 = w[2];
    w7 = w[11];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[18] = w16 + s0 + s1 + w7;
  end
  19: begin
    w15 = w[4];
    w2 = w[17];
    w16 = w[3];
    w7 = w[12];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[19] = w16 + s0 + s1 + w7;
  end
  20: begin
    w15 = w[5];
    w2 = w[18];
    w16 = w[4];
    w7 = w[13];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[20] = w16 + s0 + s1 + w7;
  end
  21: begin
    w15 = w[6];
    w2 = w[19];
    w16 = w[5];
    w7 = w[14];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[21] = w16 + s0 + s1 + w7;
  end
  22: begin
    w15 = w[7];
    w2 = w[20];
    w16 = w[6];
    w7 = w[15];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[22] = w16 + s0 + s1 + w7;
  end
  23: begin
    w15 = w[8];
    w2 = w[21];
    w16 = w[7];
    w7 = w[16];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[23] = w16 + s0 + s1 + w7;
  end
  24: begin
    w15 = w[9];
    w2 = w[22];
    w16 = w[8];
    w7 = w[17];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[24] = w16 + s0 + s1 + w7;
  end
  25: begin
    w15 = w[10];
    w2 = w[23];
    w16 = w[9];
    w7 = w[18];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[25] = w16 + s0 + s1 + w7;
  end
  26: begin
    w15 = w[11];
    w2 = w[24];
    w16 = w[10];
    w7 = w[19];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[26] = w16 + s0 + s1 + w7;
  end
  27: begin
    w15 = w[12];
    w2 = w[25];
    w16 = w[11];
    w7 = w[20];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[27] = w16 + s0 + s1 + w7;
  end
  28: begin
    w15 = w[13];
    w2 = w[26];
    w16 = w[12];
    w7 = w[21];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[28] = w16 + s0 + s1 + w7;
  end
  29: begin
    w15 = w[14];
    w2 = w[27];
    w16 = w[13];
    w7 = w[22];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[29] = w16 + s0 + s1 + w7;
  end
  30: begin
    w15 = w[15];
    w2 = w[28];
    w16 = w[14];
    w7 = w[23];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[30] = w16 + s0 + s1 + w7;
  end
  31: begin
    w15 = w[16];
    w2 = w[29];
    w16 = w[15];
    w7 = w[24];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[31] = w16 + s0 + s1 + w7;
  end
  32: begin
    w15 = w[17];
    w2 = w[30];
    w16 = w[16];
    w7 = w[25];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[32] = w16 + s0 + s1 + w7;
  end
  33: begin
    w15 = w[18];
    w2 = w[31];
    w16 = w[17];
    w7 = w[26];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[33] = w16 + s0 + s1 + w7;
  end
  34: begin
    w15 = w[19];
    w2 = w[32];
    w16 = w[18];
    w7 = w[27];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[34] = w16 + s0 + s1 + w7;
  end
  35: begin
    w15 = w[20];
    w2 = w[33];
    w16 = w[19];
    w7 = w[28];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[35] = w16 + s0 + s1 + w7;
  end
  36: begin
    w15 = w[21];
    w2 = w[34];
    w16 = w[20];
    w7 = w[29];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[36] = w16 + s0 + s1 + w7;
  end
  37: begin
    w15 = w[22];
    w2 = w[35];
    w16 = w[21];
    w7 = w[30];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[37] = w16 + s0 + s1 + w7;
  end
  38: begin
    w15 = w[23];
    w2 = w[36];
    w16 = w[22];
    w7 = w[31];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[38] = w16 + s0 + s1 + w7;
  end
  39: begin
    w15 = w[24];
    w2 = w[37];
    w16 = w[23];
    w7 = w[32];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[39] = w16 + s0 + s1 + w7;
  end
  40: begin
    w15 = w[25];
    w2 = w[38];
    w16 = w[24];
    w7 = w[33];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[40] = w16 + s0 + s1 + w7;
  end
  41: begin
    w15 = w[26];
    w2 = w[39];
    w16 = w[25];
    w7 = w[34];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[41] = w16 + s0 + s1 + w7;
  end
  42: begin
    w15 = w[27];
    w2 = w[40];
    w16 = w[26];
    w7 = w[35];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[42] = w16 + s0 + s1 + w7;
  end
  43: begin
    w15 = w[28];
    w2 = w[41];
    w16 = w[27];
    w7 = w[36];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[43] = w16 + s0 + s1 + w7;
  end
  44: begin
    w15 = w[29];
    w2 = w[42];
    w16 = w[28];
    w7 = w[37];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[44] = w16 + s0 + s1 + w7;
  end
  45: begin
    w15 = w[30];
    w2 = w[43];
    w16 = w[29];
    w7 = w[38];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[45] = w16 + s0 + s1 + w7;
  end
  46: begin
    w15 = w[31];
    w2 = w[44];
    w16 = w[30];
    w7 = w[39];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[46] = w16 + s0 + s1 + w7;
  end
  47: begin
    w15 = w[32];
    w2 = w[45];
    w16 = w[31];
    w7 = w[40];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[47] = w16 + s0 + s1 + w7;
  end
  48: begin
    w15 = w[33];
    w2 = w[46];
    w16 = w[32];
    w7 = w[41];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[48] = w16 + s0 + s1 + w7;
  end
  49: begin
    w15 = w[34];
    w2 = w[47];
    w16 = w[33];
    w7 = w[42];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[49] = w16 + s0 + s1 + w7;
  end
  50: begin
    w15 = w[35];
    w2 = w[48];
    w16 = w[34];
    w7 = w[43];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[50] = w16 + s0 + s1 + w7;
  end
  51: begin
    w15 = w[36];
    w2 = w[49];
    w16 = w[35];
    w7 = w[44];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[51] = w16 + s0 + s1 + w7;
  end
  52: begin
    w15 = w[37];
    w2 = w[50];
    w16 = w[36];
    w7 = w[45];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[52] = w16 + s0 + s1 + w7;
  end
  53: begin
    w15 = w[38];
    w2 = w[51];
    w16 = w[37];
    w7 = w[46];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[53] = w16 + s0 + s1 + w7;
  end
  54: begin
    w15 = w[39];
    w2 = w[52];
    w16 = w[38];
    w7 = w[47];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[54] = w16 + s0 + s1 + w7;
  end
  55: begin
    w15 = w[40];
    w2 = w[53];
    w16 = w[39];
    w7 = w[48];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[55] = w16 + s0 + s1 + w7;
  end
  56: begin
    w15 = w[41];
    w2 = w[54];
    w16 = w[40];
    w7 = w[49];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[56] = w16 + s0 + s1 + w7;
  end
  57: begin
    w15 = w[42];
    w2 = w[55];
    w16 = w[41];
    w7 = w[50];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[57] = w16 + s0 + s1 + w7;
  end
  58: begin
    w15 = w[43];
    w2 = w[56];
    w16 = w[42];
    w7 = w[51];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[58] = w16 + s0 + s1 + w7;
  end
  59: begin
    w15 = w[44];
    w2 = w[57];
    w16 = w[43];
    w7 = w[52];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[59] = w16 + s0 + s1 + w7;
  end
  60: begin
    w15 = w[45];
    w2 = w[58];
    w16 = w[44];
    w7 = w[53];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[60] = w16 + s0 + s1 + w7;
  end
  61: begin
    w15 = w[46];
    w2 = w[59];
    w16 = w[45];
    w7 = w[54];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[61] = w16 + s0 + s1 + w7;
  end
  62: begin
    w15 = w[47];
    w2 = w[60];
    w16 = w[46];
    w7 = w[55];
    next_state = state + 1;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[62] = w16 + s0 + s1 + w7;
  end
  63: begin
    w15 = w[48];
    w2 = w[61];
    w16 = w[47];
    w7 = w[56];
    next_state = 15;
    s0 = {w15[25:31],w15[0:24]} ^ {w15[14:31],w15[0:13]} ^ (w15 >> 3);
    s1 = {w2[15:31],w2[0:14]} ^ {w2[13:31],w2[0:12]} ^ (w2 >> 10);
    new_w[63] = w16 + s0 + s1 + w7;
  end
  endcase
  if(msa_en == 1) begin
      next_state = 16;
      new_w[0:15] = chunk;
  end
  end
endmodule