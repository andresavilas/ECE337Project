// $Id: $
// File name:   miner_core_comp.sv
// Created:     4/20/2015
// Author:      Andres Avila
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Compression Function
module miner_core_comp (
  input wire comp_en,
  input wire clk,
  input wire n_rst,
  input wire [0:63] [0:31] w,
  input wire [0:7] [0:31] first_h,
  output logic [0:7] [0:31] h
);
  reg [0:6] state;
  reg [0:6] next_state;
  reg [0:31] S1;
  reg [0:31] S0;
  reg [0:31] temp1;
  reg [0:31] temp2;
  reg [0:31] maj;
  reg [0:31] ch;
  logic [0:7] [0:31] new_h;
  wire [0:63] [0:31] k = {32'h428a2f98, 32'h71374491, 32'hb5c0fbcf, 32'he9b5dba5, 32'h3956c25b, 32'h59f111f1, 32'h923f82a4, 32'hab1c5ed5, 32'hd807aa98, 32'h12835b01, 32'h243185be, 32'h550c7dc3, 32'h72be5d74, 32'h80deb1fe, 32'h9bdc06a7, 32'hc19bf174,
   32'he49b69c1, 32'hefbe4786, 32'h0fc19dc6, 32'h240ca1cc, 32'h2de92c6f, 32'h4a7484aa, 32'h5cb0a9dc, 32'h76f988da,
   32'h983e5152, 32'ha831c66d, 32'hb00327c8, 32'hbf597fc7, 32'hc6e00bf3, 32'hd5a79147, 32'h06ca6351, 32'h14292967,
   32'h27b70a85, 32'h2e1b2138, 32'h4d2c6dfc, 32'h53380d13, 32'h650a7354, 32'h766a0abb, 32'h81c2c92e, 32'h92722c85,
   32'ha2bfe8a1, 32'ha81a664b, 32'hc24b8b70, 32'hc76c51a3, 32'hd192e819, 32'hd6990624, 32'hf40e3585, 32'h106aa070,
   32'h19a4c116, 32'h1e376c08, 32'h2748774c, 32'h34b0bcb5, 32'h391c0cb3, 32'h4ed8aa4a, 32'h5b9cca4f, 32'h682e6ff3,
   32'h748f82ee, 32'h78a5636f, 32'h84c87814, 32'h8cc70208, 32'h90befffa, 32'ha4506ceb, 32'hbef9a3f7, 32'hc67178f2};
  always_ff @ (posedge clk, negedge n_rst) begin
    if(n_rst == 0) begin
      h <= 0;
      state <= 0;
    end else begin
      h <= new_h;
      state <= next_state;
    end
  end
  always_comb begin
    next_state = state;
    new_h = h;
    case (state)
      0: begin
        if(comp_en == 1) begin
          next_state = 1;
          S1 = {first_h[4][26:31],first_h[4][0:25]} ^ {first_h[4][21:31],first_h[4][0:20]} ^ {first_h[4][7:31],first_h[4][0:6]};
          ch = (first_h[4] & first_h[5]) ^ ((~first_h[4]) & first_h[6]);
          temp1 = first_h[7] + S1 + ch + k[0] + w[0];
          S0 = {first_h[0][30:31],first_h[0][0:29]} ^ {first_h[0][19:31],first_h[0][0:18]} ^ {first_h[0][10:31],first_h[0][0:9]}; 
          maj = (first_h[0] & first_h[1]) ^ (first_h[0] & first_h[2]) ^ {first_h[1] & first_h[2]};
          temp2 = S0 + maj;
          new_h[0] = temp1 + temp2;
          new_h[1] = first_h[0];
          new_h[2] = first_h[1];
          new_h[3] = first_h[2];
          new_h[4] = first_h[3] + temp1;
          new_h[5] = first_h[4];
          new_h[6] = first_h[5];
          new_h[7] = first_h[6];  
        end
      end
       1: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[1] + w[1];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  2: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[2] + w[2];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  3: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[3] + w[3];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  4: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[4] + w[4];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  5: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[5] + w[5];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  6: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[6] + w[6];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  7: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[7] + w[7];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  8: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[8] + w[8];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  9: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[9] + w[9];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  10: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[10] + w[10];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  11: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[11] + w[11];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  12: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[12] + w[12];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  13: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[13] + w[13];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  14: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[14] + w[14];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  15: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[15] + w[15];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  16: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[16] + w[16];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  17: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[17] + w[17];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  18: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[18] + w[18];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  19: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[19] + w[19];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  20: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[20] + w[20];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  21: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[21] + w[21];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  22: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[22] + w[22];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  23: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[23] + w[23];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  24: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[24] + w[24];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  25: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[25] + w[25];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  26: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[26] + w[26];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  27: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[27] + w[27];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  28: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[28] + w[28];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  29: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[29] + w[29];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  30: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[30] + w[30];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  31: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[31] + w[31];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  32: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[32] + w[32];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  33: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[33] + w[33];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  34: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[34] + w[34];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  35: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[35] + w[35];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  36: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[36] + w[36];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  37: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[37] + w[37];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  38: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[38] + w[38];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  39: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[39] + w[39];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  40: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[40] + w[40];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  41: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[41] + w[41];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  42: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[42] + w[42];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  43: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[43] + w[43];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  44: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[44] + w[44];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  45: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[45] + w[45];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  46: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[46] + w[46];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  47: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[47] + w[47];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  48: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[48] + w[48];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  49: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[49] + w[49];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  50: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[50] + w[50];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  51: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[51] + w[51];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  52: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[52] + w[52];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  53: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[53] + w[53];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  54: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[54] + w[54];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  55: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[55] + w[55];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  56: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[56] + w[56];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  57: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[57] + w[57];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  58: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[58] + w[58];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  59: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[59] + w[59];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  60: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[60] + w[60];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  61: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[61] + w[61];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  62: begin
    next_state = state + 1;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[62] + w[62];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
  63: begin
    next_state = 0;
    S1 = {h[4][26:31],h[4][0:25]} ^ {h[4][21:31],h[4][0:20]} ^ {h[4][7:31],h[4][0:6]};
    ch = (h[4] & h[5]) ^ ((~h[4]) & h[6]);
    temp1 = h[7] + S1 + ch + k[63] + w[63];
    S0 = {h[0][30:31],h[0][0:29]} ^ {h[0][19:31],h[0][0:18]} ^ {h[0][10:31],h[0][0:9]};
    maj = (h[0] & h[1]) ^ (h[0] & h[2]) ^ {h[1] & h[2]};
    temp2 = S0 + maj;
    new_h[0] = temp1 + temp2;
    new_h[1] = h[0];
    new_h[2] = h[1];
    new_h[3] = h[2];
    new_h[4] = h[3] + temp1;
    new_h[5] = h[4];
    new_h[6] = h[5];
    new_h[7] = h[6];
  end
endcase
  end    
endmodule 