library verilog;
use verilog.vl_types.all;
entity tb_uartrx_sv_unit is
end tb_uartrx_sv_unit;
