library verilog;
use verilog.vl_types.all;
entity tb_uart_tx_sv_unit is
end tb_uart_tx_sv_unit;
