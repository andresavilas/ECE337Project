library verilog;
use verilog.vl_types.all;
entity tb_uartrx is
end tb_uartrx;
